---------------------------------------------------------------------
-- TITLE: Random Access Memory for Xilinx
-- AUTHOR: Steve Rhoads (rhoadss@yahoo.com)
-- DATE CREATED: 11/06/05
-- FILENAME: cache_ram.vhd
-- PROJECT: Plasma CPU core
-- COPYRIGHT: Software placed into the public domain by the author.
--    Software 'as is' without warranty.  Author liable for nothing.
-- DESCRIPTION:
--    Implements Plasma Cache RAM as RAMB 
--    The file is configurable up to 64KB, in blocks of 8 KB.
--    The Cache Data RAM uses only the lower 4KB of block0
--
-- MEMORY MAP
--    0000..1FFF : 8KB   8KB  block0
--    2000..3FFF : 8KB  16KB  block1 
--    4000..5FFF : 8KB  24KB  block2
--    6000..7FFF : 8KB  32KB  block3
--    8000..9FFF : 8KB  40KB  block4
--    A000..BFFF : 8KB  48KB  block5
--    C000..DFFF : 8KB  56KB  block6
--    E000..FFFF : 8KB  64KB  block7
---------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use work.mlite_pack.all;

library UNISIM;
use UNISIM.vcomponents.all;

entity cache_ram is
   generic( block_count : integer := 1); 
   port(clk               : in std_logic;
        enable            : in std_logic;
        write_byte_enable : in std_logic_vector(3 downto 0);
        address           : in std_logic_vector(31 downto 2);
        data_write        : in std_logic_vector(31 downto 0);
        data_read         : out std_logic_vector(31 downto 0));
end; --entity ram

architecture logic of cache_ram is
   --type
   --type mem32_vector IS ARRAY (NATURAL RANGE<>) OF std_logic_vector(31 downto 0);

   --Which 8KB block
   --alias block_sel: std_logic_vector(2 downto 0) is address(15 downto 13);

   --Address within a 8KB block (without lower two bits)
   alias block_addr : std_logic_vector(10 downto 0) is address(12 downto 2);

   --Block enable with 1 bit per memory block
   --signal block_enable: std_logic_vector(7 downto 0);

   --Block Data Out
   --signal block_do: mem32_vector(7 downto 0);

   --Remember which block was selected
   --signal block_sel_buf: std_logic_vector(2 downto 0);

begin
   -- block_enable<= "00000001" when (enable='1') and (block_sel="000") else 
                  -- "00000010" when (enable='1') and (block_sel="001") else 
                  -- "00000100" when (enable='1') and (block_sel="010") else 
                  -- "00001000" when (enable='1') and (block_sel="011") else 
                  -- "00010000" when (enable='1') and (block_sel="100") else 
                  -- "00100000" when (enable='1') and (block_sel="101") else 
                  -- "01000000" when (enable='1') and (block_sel="110") else 
                  -- "10000000" when (enable='1') and (block_sel="111") else
                  -- "00000000";
  
   -- proc_blocksel: process (clk, block_sel) is
   -- begin
      -- if rising_edge(clk) then 
         -- block_sel_buf <= block_sel;
      -- end if;
   -- end process;

   -- proc_do: process (block_do, block_sel_buf) is
   -- begin
      -- data_read <= block_do(conv_integer(block_sel_buf));
   -- end process;
	
	-- BLOCKS generation
   block0: if (block_count > 0) generate
	begin

    ram_byte3 : RAMB16_S9
   generic map (
INIT_00 => X"000000000000000000000000000000000000000000000000000000000c080400",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
)
    port map (
      DO   => data_read(31 downto 24), 
      DOP  => open, 
      ADDR => block_addr,
      CLK  => clk, 
      DI   => data_write(31 downto 24),
      DIP  => ZERO(0 downto 0),
      EN   => enable,
      SSR  => ZERO(0),
      WE   => write_byte_enable(3));

    ram_byte2 : RAMB16_S9
   generic map (
INIT_00 => X"000000000000000000000000000000000000000000000000000000000d090501",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
)
    port map (
      DO   => data_read(23 downto 16),
      DOP  => open, 
      ADDR => block_addr,
      CLK  => clk, 
      DI   => data_write(23 downto 16),
      DIP  => ZERO(0 downto 0),
      EN   => enable,
      SSR  => ZERO(0),
      WE   => write_byte_enable(2));
	
    ram_byte1 : RAMB16_S9
   generic map (
INIT_00 => X"000000000000000000000000000000000000000000000000000000000e0a0602",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
)
    port map (
      DO   => data_read(15 downto 8),
      DOP  => open, 
      ADDR => block_addr,
      CLK  => clk, 
      DI   => data_write(15 downto 8),
      DIP  => ZERO(0 downto 0),
      EN   => enable,
      SSR  => ZERO(0),
      WE   => write_byte_enable(1));

    ram_byte0 : RAMB16_S9
   generic map (
INIT_00 => X"000000000000000000000000000000000000000000000000000000000f0b0703",
INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
)
    port map (
      DO   => data_read(7 downto 0),
      DOP  => open, 
      ADDR => block_addr,
      CLK  => clk, 
      DI   => data_write(7 downto 0),
      DIP  => ZERO(0 downto 0),
      EN   => enable,
      SSR  => ZERO(0),
      WE   => write_byte_enable(0));
   end generate; --block0
	

   -- block1: if (block_count > 1) generate
	-- begin

    -- ram_byte3 : RAMB16_S9
   -- generic map (
-- INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
-- )
    -- port map (
      -- DO   => block_do(1)(31 downto 24), 
      -- DOP  => open, 
      -- ADDR => block_addr,
      -- CLK  => clk, 
      -- DI   => data_write(31 downto 24),
      -- DIP  => ZERO(0 downto 0),
      -- EN   => block_enable(1),
      -- SSR  => ZERO(0),
      -- WE   => write_byte_enable(3));

    -- ram_byte2 : RAMB16_S9
   -- generic map (
-- INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
-- )
    -- port map (
      -- DO   => block_do(1)(23 downto 16),
      -- DOP  => open, 
      -- ADDR => block_addr,
      -- CLK  => clk, 
      -- DI   => data_write(23 downto 16),
      -- DIP  => ZERO(0 downto 0),
      -- EN   => block_enable(1),
      -- SSR  => ZERO(0),
      -- WE   => write_byte_enable(2));
	
    -- ram_byte1 : RAMB16_S9
   -- generic map (
-- INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
-- )
    -- port map (
      -- DO   => block_do(1)(15 downto 8),
      -- DOP  => open, 
      -- ADDR => block_addr,
      -- CLK  => clk, 
      -- DI   => data_write(15 downto 8),
      -- DIP  => ZERO(0 downto 0),
      -- EN   => block_enable(1),
      -- SSR  => ZERO(0),
      -- WE   => write_byte_enable(1));

    -- ram_byte0 : RAMB16_S9
   -- generic map (
-- INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
-- )
    -- port map (
      -- DO   => block_do(1)(7 downto 0),
      -- DOP  => open, 
      -- ADDR => block_addr,
      -- CLK  => clk, 
      -- DI   => data_write(7 downto 0),
      -- DIP  => ZERO(0 downto 0),
      -- EN   => block_enable(1),
      -- SSR  => ZERO(0),
      -- WE   => write_byte_enable(0));
		
   -- end generate; --block1
	

   -- block2: if (block_count > 2) generate
	-- begin

    -- ram_byte3 : RAMB16_S9
   -- generic map (
-- INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
-- )
    -- port map (
      -- DO   => block_do(2)(31 downto 24), 
      -- DOP  => open, 
      -- ADDR => block_addr,
      -- CLK  => clk, 
      -- DI   => data_write(31 downto 24),
      -- DIP  => ZERO(0 downto 0),
      -- EN   => block_enable(2),
      -- SSR  => ZERO(0),
      -- WE   => write_byte_enable(3));

    -- ram_byte2 : RAMB16_S9
   -- generic map (
-- INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
-- )
    -- port map (
      -- DO   => block_do(2)(23 downto 16),
      -- DOP  => open, 
      -- ADDR => block_addr,
      -- CLK  => clk, 
      -- DI   => data_write(23 downto 16),
      -- DIP  => ZERO(0 downto 0),
      -- EN   => block_enable(2),
      -- SSR  => ZERO(0),
      -- WE   => write_byte_enable(2));
	
    -- ram_byte1 : RAMB16_S9
   -- generic map (
-- INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
-- )
    -- port map (
      -- DO   => block_do(2)(15 downto 8),
      -- DOP  => open, 
      -- ADDR => block_addr,
      -- CLK  => clk, 
      -- DI   => data_write(15 downto 8),
      -- DIP  => ZERO(0 downto 0),
      -- EN   => block_enable(2),
      -- SSR  => ZERO(0),
      -- WE   => write_byte_enable(1));

    -- ram_byte0 : RAMB16_S9
   -- generic map (
-- INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
-- )
    -- port map (
      -- DO   => block_do(2)(7 downto 0),
      -- DOP  => open, 
      -- ADDR => block_addr,
      -- CLK  => clk, 
      -- DI   => data_write(7 downto 0),
      -- DIP  => ZERO(0 downto 0),
      -- EN   => block_enable(2),
      -- SSR  => ZERO(0),
      -- WE   => write_byte_enable(0));
		
   -- end generate; --block2


   -- block3: if (block_count > 3) generate
	-- begin

    -- ram_byte3 : RAMB16_S9
   -- generic map (
-- INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
-- )
    -- port map (
      -- DO   => block_do(3)(31 downto 24), 
      -- DOP  => open, 
      -- ADDR => block_addr,
      -- CLK  => clk, 
      -- DI   => data_write(31 downto 24),
      -- DIP  => ZERO(0 downto 0),
      -- EN   => block_enable(3),
      -- SSR  => ZERO(0),
      -- WE   => write_byte_enable(3));

    -- ram_byte2 : RAMB16_S9
   -- generic map (
-- INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
-- )
    -- port map (
      -- DO   => block_do(3)(23 downto 16),
      -- DOP  => open, 
      -- ADDR => block_addr,
      -- CLK  => clk, 
      -- DI   => data_write(23 downto 16),
      -- DIP  => ZERO(0 downto 0),
      -- EN   => block_enable(3),
      -- SSR  => ZERO(0),
      -- WE   => write_byte_enable(2));
	
    -- ram_byte1 : RAMB16_S9
   -- generic map (
-- INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
-- )
    -- port map (
      -- DO   => block_do(3)(15 downto 8),
      -- DOP  => open, 
      -- ADDR => block_addr,
      -- CLK  => clk, 
      -- DI   => data_write(15 downto 8),
      -- DIP  => ZERO(0 downto 0),
      -- EN   => block_enable(3),
      -- SSR  => ZERO(0),
      -- WE   => write_byte_enable(1));

    -- ram_byte0 : RAMB16_S9
   -- generic map (
-- INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
-- )
    -- port map (
      -- DO   => block_do(3)(7 downto 0),
      -- DOP  => open, 
      -- ADDR => block_addr,
      -- CLK  => clk, 
      -- DI   => data_write(7 downto 0),
      -- DIP  => ZERO(0 downto 0),
      -- EN   => block_enable(3),
      -- SSR  => ZERO(0),
      -- WE   => write_byte_enable(0));
		
   -- end generate; --block3


   -- block4: if (block_count > 4) generate
	-- begin

    -- ram_byte3 : RAMB16_S9
   -- generic map (
-- INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
-- )
    -- port map (
      -- DO   => block_do(4)(31 downto 24), 
      -- DOP  => open, 
      -- ADDR => block_addr,
      -- CLK  => clk, 
      -- DI   => data_write(31 downto 24),
      -- DIP  => ZERO(0 downto 0),
      -- EN   => block_enable(4),
      -- SSR  => ZERO(0),
      -- WE   => write_byte_enable(3));

    -- ram_byte2 : RAMB16_S9
   -- generic map (
-- INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
-- )
    -- port map (
      -- DO   => block_do(4)(23 downto 16),
      -- DOP  => open, 
      -- ADDR => block_addr,
      -- CLK  => clk, 
      -- DI   => data_write(23 downto 16),
      -- DIP  => ZERO(0 downto 0),
      -- EN   => block_enable(4),
      -- SSR  => ZERO(0),
      -- WE   => write_byte_enable(2));
	
    -- ram_byte1 : RAMB16_S9
   -- generic map (
-- INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
-- )
    -- port map (
      -- DO   => block_do(4)(15 downto 8),
      -- DOP  => open, 
      -- ADDR => block_addr,
      -- CLK  => clk, 
      -- DI   => data_write(15 downto 8),
      -- DIP  => ZERO(0 downto 0),
      -- EN   => block_enable(4),
      -- SSR  => ZERO(0),
      -- WE   => write_byte_enable(1));

    -- ram_byte0 : RAMB16_S9
   -- generic map (
-- INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
-- )
    -- port map (
      -- DO   => block_do(4)(7 downto 0),
      -- DOP  => open, 
      -- ADDR => block_addr,
      -- CLK  => clk, 
      -- DI   => data_write(7 downto 0),
      -- DIP  => ZERO(0 downto 0),
      -- EN   => block_enable(4),
      -- SSR  => ZERO(0),
      -- WE   => write_byte_enable(0));
		
   -- end generate; --block4


   -- block5: if (block_count > 5) generate
	-- begin

    -- ram_byte3 : RAMB16_S9
   -- generic map (
-- INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
-- )
    -- port map (
      -- DO   => block_do(5)(31 downto 24), 
      -- DOP  => open, 
      -- ADDR => block_addr,
      -- CLK  => clk, 
      -- DI   => data_write(31 downto 24),
      -- DIP  => ZERO(0 downto 0),
      -- EN   => block_enable(5),
      -- SSR  => ZERO(0),
      -- WE   => write_byte_enable(3));

    -- ram_byte2 : RAMB16_S9
   -- generic map (
-- INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
-- )
    -- port map (
      -- DO   => block_do(5)(23 downto 16),
      -- DOP  => open, 
      -- ADDR => block_addr,
      -- CLK  => clk, 
      -- DI   => data_write(23 downto 16),
      -- DIP  => ZERO(0 downto 0),
      -- EN   => block_enable(5),
      -- SSR  => ZERO(0),
      -- WE   => write_byte_enable(2));
	
    -- ram_byte1 : RAMB16_S9
   -- generic map (
-- INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
-- )
    -- port map (
      -- DO   => block_do(5)(15 downto 8),
      -- DOP  => open, 
      -- ADDR => block_addr,
      -- CLK  => clk, 
      -- DI   => data_write(15 downto 8),
      -- DIP  => ZERO(0 downto 0),
      -- EN   => block_enable(5),
      -- SSR  => ZERO(0),
      -- WE   => write_byte_enable(1));

    -- ram_byte0 : RAMB16_S9
   -- generic map (
-- INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
-- )
    -- port map (
      -- DO   => block_do(5)(7 downto 0),
      -- DOP  => open, 
      -- ADDR => block_addr,
      -- CLK  => clk, 
      -- DI   => data_write(7 downto 0),
      -- DIP  => ZERO(0 downto 0),
      -- EN   => block_enable(5),
      -- SSR  => ZERO(0),
      -- WE   => write_byte_enable(0));
		
   -- end generate; --block5


   -- block6: if (block_count > 6) generate
	-- begin

    -- ram_byte3 : RAMB16_S9
   -- generic map (
-- INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
-- )
    -- port map (
      -- DO   => block_do(6)(31 downto 24), 
      -- DOP  => open, 
      -- ADDR => block_addr,
      -- CLK  => clk, 
      -- DI   => data_write(31 downto 24),
      -- DIP  => ZERO(0 downto 0),
      -- EN   => block_enable(6),
      -- SSR  => ZERO(0),
      -- WE   => write_byte_enable(3));

    -- ram_byte2 : RAMB16_S9
   -- generic map (
-- INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
-- )
    -- port map (
      -- DO   => block_do(6)(23 downto 16),
      -- DOP  => open, 
      -- ADDR => block_addr,
      -- CLK  => clk, 
      -- DI   => data_write(23 downto 16),
      -- DIP  => ZERO(0 downto 0),
      -- EN   => block_enable(6),
      -- SSR  => ZERO(0),
      -- WE   => write_byte_enable(2));
	
    -- ram_byte1 : RAMB16_S9
   -- generic map (
-- INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
-- )
    -- port map (
      -- DO   => block_do(6)(15 downto 8),
      -- DOP  => open, 
      -- ADDR => block_addr,
      -- CLK  => clk, 
      -- DI   => data_write(15 downto 8),
      -- DIP  => ZERO(0 downto 0),
      -- EN   => block_enable(6),
      -- SSR  => ZERO(0),
      -- WE   => write_byte_enable(1));

    -- ram_byte0 : RAMB16_S9
   -- generic map (
-- INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
-- )
    -- port map (
      -- DO   => block_do(6)(7 downto 0),
      -- DOP  => open, 
      -- ADDR => block_addr,
      -- CLK  => clk, 
      -- DI   => data_write(7 downto 0),
      -- DIP  => ZERO(0 downto 0),
      -- EN   => block_enable(6),
      -- SSR  => ZERO(0),
      -- WE   => write_byte_enable(0));
		
   -- end generate; --block6


   -- block7: if (block_count > 7) generate
	-- begin

    -- ram_byte3 : RAMB16_S9
   -- generic map (
-- INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
-- )
    -- port map (
      -- DO   => block_do(7)(31 downto 24), 
      -- DOP  => open, 
      -- ADDR => block_addr,
      -- CLK  => clk, 
      -- DI   => data_write(31 downto 24),
      -- DIP  => ZERO(0 downto 0),
      -- EN   => block_enable(7),
      -- SSR  => ZERO(0),
      -- WE   => write_byte_enable(3));

    -- ram_byte2 : RAMB16_S9
   -- generic map (
-- INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
-- )
    -- port map (
      -- DO   => block_do(7)(23 downto 16),
      -- DOP  => open, 
      -- ADDR => block_addr,
      -- CLK  => clk, 
      -- DI   => data_write(23 downto 16),
      -- DIP  => ZERO(0 downto 0),
      -- EN   => block_enable(7),
      -- SSR  => ZERO(0),
      -- WE   => write_byte_enable(2));
	
    -- ram_byte1 : RAMB16_S9
   -- generic map (
-- INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
-- )
    -- port map (
      -- DO   => block_do(7)(15 downto 8),
      -- DOP  => open, 
      -- ADDR => block_addr,
      -- CLK  => clk, 
      -- DI   => data_write(15 downto 8),
      -- DIP  => ZERO(0 downto 0),
      -- EN   => block_enable(7),
      -- SSR  => ZERO(0),
      -- WE   => write_byte_enable(1));

    -- ram_byte0 : RAMB16_S9
   -- generic map (
-- INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
-- INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000"
-- )
    -- port map (
      -- DO   => block_do(7)(7 downto 0),
      -- DOP  => open, 
      -- ADDR => block_addr,
      -- CLK  => clk, 
      -- DI   => data_write(7 downto 0),
      -- DIP  => ZERO(0 downto 0),
      -- EN   => block_enable(7),
      -- SSR  => ZERO(0),
      -- WE   => write_byte_enable(0));
		
   -- end generate; --block7

end; --architecture logic
