library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use IEEE.std_logic_arith.all;

entity CSA is
port(
in1 : in std_logic_vector(31 downto 0);
in2 : in std_logic_vector(31 downto 0);
out1 : out std_logic_vector(62 downto 0);
out2 : out std_logic_vector(62 downto 0));
end;

architecture structural of CSA is

	component FA is
	port(in1 : in std_logic;
		in2 : in std_logic;
		c_in : in std_logic;
		sum : out std_logic;
		c_out : out std_logic);
	end component;

--signals for iteration 0
signal CSA_sum_0_2_0, CSA_carry_0_2_0, CSA_sum_0_3_0, CSA_carry_0_3_0, CSA_sum_0_4_0, CSA_carry_0_4_0, CSA_sum_0_5_0, CSA_carry_0_5_0, CSA_sum_0_5_1, CSA_carry_0_5_1, CSA_sum_0_6_0, CSA_carry_0_6_0, CSA_sum_0_6_1, CSA_carry_0_6_1, CSA_sum_0_7_0, CSA_carry_0_7_0, CSA_sum_0_7_1, CSA_carry_0_7_1, CSA_sum_0_8_0, CSA_carry_0_8_0, CSA_sum_0_8_1, CSA_carry_0_8_1, CSA_sum_0_8_2, CSA_carry_0_8_2, CSA_sum_0_9_0, CSA_carry_0_9_0, CSA_sum_0_9_1, CSA_carry_0_9_1, CSA_sum_0_9_2, CSA_carry_0_9_2, CSA_sum_0_10_0, CSA_carry_0_10_0, CSA_sum_0_10_1, CSA_carry_0_10_1, CSA_sum_0_10_2, CSA_carry_0_10_2, CSA_sum_0_11_0, CSA_carry_0_11_0, CSA_sum_0_11_1, CSA_carry_0_11_1, CSA_sum_0_11_2, CSA_carry_0_11_2, CSA_sum_0_11_3, CSA_carry_0_11_3, CSA_sum_0_12_0, CSA_carry_0_12_0, CSA_sum_0_12_1, CSA_carry_0_12_1, CSA_sum_0_12_2, CSA_carry_0_12_2, CSA_sum_0_12_3, CSA_carry_0_12_3, CSA_sum_0_13_0, CSA_carry_0_13_0, CSA_sum_0_13_1, CSA_carry_0_13_1, CSA_sum_0_13_2, CSA_carry_0_13_2, CSA_sum_0_13_3, CSA_carry_0_13_3, CSA_sum_0_14_0, CSA_carry_0_14_0, CSA_sum_0_14_1, CSA_carry_0_14_1, CSA_sum_0_14_2, CSA_carry_0_14_2, CSA_sum_0_14_3, CSA_carry_0_14_3, CSA_sum_0_14_4, CSA_carry_0_14_4, CSA_sum_0_15_0, CSA_carry_0_15_0, CSA_sum_0_15_1, CSA_carry_0_15_1, CSA_sum_0_15_2, CSA_carry_0_15_2, CSA_sum_0_15_3, CSA_carry_0_15_3, CSA_sum_0_15_4, CSA_carry_0_15_4, CSA_sum_0_16_0, CSA_carry_0_16_0, CSA_sum_0_16_1, CSA_carry_0_16_1, CSA_sum_0_16_2, CSA_carry_0_16_2, CSA_sum_0_16_3, CSA_carry_0_16_3, CSA_sum_0_16_4, CSA_carry_0_16_4, CSA_sum_0_17_0, CSA_carry_0_17_0, CSA_sum_0_17_1, CSA_carry_0_17_1, CSA_sum_0_17_2, CSA_carry_0_17_2, CSA_sum_0_17_3, CSA_carry_0_17_3, CSA_sum_0_17_4, CSA_carry_0_17_4, CSA_sum_0_17_5, CSA_carry_0_17_5, CSA_sum_0_18_0, CSA_carry_0_18_0, CSA_sum_0_18_1, CSA_carry_0_18_1, CSA_sum_0_18_2, CSA_carry_0_18_2, CSA_sum_0_18_3, CSA_carry_0_18_3, CSA_sum_0_18_4, CSA_carry_0_18_4, CSA_sum_0_18_5, CSA_carry_0_18_5, CSA_sum_0_19_0, CSA_carry_0_19_0, CSA_sum_0_19_1, CSA_carry_0_19_1, CSA_sum_0_19_2, CSA_carry_0_19_2, CSA_sum_0_19_3, CSA_carry_0_19_3, CSA_sum_0_19_4, CSA_carry_0_19_4, CSA_sum_0_19_5, CSA_carry_0_19_5, CSA_sum_0_20_0, CSA_carry_0_20_0, CSA_sum_0_20_1, CSA_carry_0_20_1, CSA_sum_0_20_2, CSA_carry_0_20_2, CSA_sum_0_20_3, CSA_carry_0_20_3, CSA_sum_0_20_4, CSA_carry_0_20_4, CSA_sum_0_20_5, CSA_carry_0_20_5, CSA_sum_0_20_6, CSA_carry_0_20_6, CSA_sum_0_21_0, CSA_carry_0_21_0, CSA_sum_0_21_1, CSA_carry_0_21_1, CSA_sum_0_21_2, CSA_carry_0_21_2, CSA_sum_0_21_3, CSA_carry_0_21_3, CSA_sum_0_21_4, CSA_carry_0_21_4, CSA_sum_0_21_5, CSA_carry_0_21_5, CSA_sum_0_21_6, CSA_carry_0_21_6, CSA_sum_0_22_0, CSA_carry_0_22_0, CSA_sum_0_22_1, CSA_carry_0_22_1, CSA_sum_0_22_2, CSA_carry_0_22_2, CSA_sum_0_22_3, CSA_carry_0_22_3, CSA_sum_0_22_4, CSA_carry_0_22_4, CSA_sum_0_22_5, CSA_carry_0_22_5, CSA_sum_0_22_6, CSA_carry_0_22_6, CSA_sum_0_23_0, CSA_carry_0_23_0, CSA_sum_0_23_1, CSA_carry_0_23_1, CSA_sum_0_23_2, CSA_carry_0_23_2, CSA_sum_0_23_3, CSA_carry_0_23_3, CSA_sum_0_23_4, CSA_carry_0_23_4, CSA_sum_0_23_5, CSA_carry_0_23_5, CSA_sum_0_23_6, CSA_carry_0_23_6, CSA_sum_0_23_7, CSA_carry_0_23_7, CSA_sum_0_24_0, CSA_carry_0_24_0, CSA_sum_0_24_1, CSA_carry_0_24_1, CSA_sum_0_24_2, CSA_carry_0_24_2, CSA_sum_0_24_3, CSA_carry_0_24_3, CSA_sum_0_24_4, CSA_carry_0_24_4, CSA_sum_0_24_5, CSA_carry_0_24_5, CSA_sum_0_24_6, CSA_carry_0_24_6, CSA_sum_0_24_7, CSA_carry_0_24_7, CSA_sum_0_25_0, CSA_carry_0_25_0, CSA_sum_0_25_1, CSA_carry_0_25_1, CSA_sum_0_25_2, CSA_carry_0_25_2, CSA_sum_0_25_3, CSA_carry_0_25_3, CSA_sum_0_25_4, CSA_carry_0_25_4, CSA_sum_0_25_5, CSA_carry_0_25_5, CSA_sum_0_25_6, CSA_carry_0_25_6, CSA_sum_0_25_7, CSA_carry_0_25_7, CSA_sum_0_26_0, CSA_carry_0_26_0, CSA_sum_0_26_1, CSA_carry_0_26_1, CSA_sum_0_26_2, CSA_carry_0_26_2, CSA_sum_0_26_3, CSA_carry_0_26_3, CSA_sum_0_26_4, CSA_carry_0_26_4, CSA_sum_0_26_5, CSA_carry_0_26_5, CSA_sum_0_26_6, CSA_carry_0_26_6, CSA_sum_0_26_7, CSA_carry_0_26_7, CSA_sum_0_26_8, CSA_carry_0_26_8, CSA_sum_0_27_0, CSA_carry_0_27_0, CSA_sum_0_27_1, CSA_carry_0_27_1, CSA_sum_0_27_2, CSA_carry_0_27_2, CSA_sum_0_27_3, CSA_carry_0_27_3, CSA_sum_0_27_4, CSA_carry_0_27_4, CSA_sum_0_27_5, CSA_carry_0_27_5, CSA_sum_0_27_6, CSA_carry_0_27_6, CSA_sum_0_27_7, CSA_carry_0_27_7, CSA_sum_0_27_8, CSA_carry_0_27_8, CSA_sum_0_28_0, CSA_carry_0_28_0, CSA_sum_0_28_1, CSA_carry_0_28_1, CSA_sum_0_28_2, CSA_carry_0_28_2, CSA_sum_0_28_3, CSA_carry_0_28_3, CSA_sum_0_28_4, CSA_carry_0_28_4, CSA_sum_0_28_5, CSA_carry_0_28_5, CSA_sum_0_28_6, CSA_carry_0_28_6, CSA_sum_0_28_7, CSA_carry_0_28_7, CSA_sum_0_28_8, CSA_carry_0_28_8, CSA_sum_0_29_0, CSA_carry_0_29_0, CSA_sum_0_29_1, CSA_carry_0_29_1, CSA_sum_0_29_2, CSA_carry_0_29_2, CSA_sum_0_29_3, CSA_carry_0_29_3, CSA_sum_0_29_4, CSA_carry_0_29_4, CSA_sum_0_29_5, CSA_carry_0_29_5, CSA_sum_0_29_6, CSA_carry_0_29_6, CSA_sum_0_29_7, CSA_carry_0_29_7, CSA_sum_0_29_8, CSA_carry_0_29_8, CSA_sum_0_29_9, CSA_carry_0_29_9, CSA_sum_0_30_0, CSA_carry_0_30_0, CSA_sum_0_30_1, CSA_carry_0_30_1, CSA_sum_0_30_2, CSA_carry_0_30_2, CSA_sum_0_30_3, CSA_carry_0_30_3, CSA_sum_0_30_4, CSA_carry_0_30_4, CSA_sum_0_30_5, CSA_carry_0_30_5, CSA_sum_0_30_6, CSA_carry_0_30_6, CSA_sum_0_30_7, CSA_carry_0_30_7, CSA_sum_0_30_8, CSA_carry_0_30_8, CSA_sum_0_30_9, CSA_carry_0_30_9, CSA_sum_0_31_0, CSA_carry_0_31_0, CSA_sum_0_31_1, CSA_carry_0_31_1, CSA_sum_0_31_2, CSA_carry_0_31_2, CSA_sum_0_31_3, CSA_carry_0_31_3, CSA_sum_0_31_4, CSA_carry_0_31_4, CSA_sum_0_31_5, CSA_carry_0_31_5, CSA_sum_0_31_6, CSA_carry_0_31_6, CSA_sum_0_31_7, CSA_carry_0_31_7, CSA_sum_0_31_8, CSA_carry_0_31_8, CSA_sum_0_31_9, CSA_carry_0_31_9, CSA_sum_0_32_0, CSA_carry_0_32_0, CSA_sum_0_32_1, CSA_carry_0_32_1, CSA_sum_0_32_2, CSA_carry_0_32_2, CSA_sum_0_32_3, CSA_carry_0_32_3, CSA_sum_0_32_4, CSA_carry_0_32_4, CSA_sum_0_32_5, CSA_carry_0_32_5, CSA_sum_0_32_6, CSA_carry_0_32_6, CSA_sum_0_32_7, CSA_carry_0_32_7, CSA_sum_0_32_8, CSA_carry_0_32_8, CSA_sum_0_32_9, CSA_carry_0_32_9, CSA_sum_0_33_0, CSA_carry_0_33_0, CSA_sum_0_33_1, CSA_carry_0_33_1, CSA_sum_0_33_2, CSA_carry_0_33_2, CSA_sum_0_33_3, CSA_carry_0_33_3, CSA_sum_0_33_4, CSA_carry_0_33_4, CSA_sum_0_33_5, CSA_carry_0_33_5, CSA_sum_0_33_6, CSA_carry_0_33_6, CSA_sum_0_33_7, CSA_carry_0_33_7, CSA_sum_0_33_8, CSA_carry_0_33_8, CSA_sum_0_33_9, CSA_carry_0_33_9, CSA_sum_0_34_0, CSA_carry_0_34_0, CSA_sum_0_34_1, CSA_carry_0_34_1, CSA_sum_0_34_2, CSA_carry_0_34_2, CSA_sum_0_34_3, CSA_carry_0_34_3, CSA_sum_0_34_4, CSA_carry_0_34_4, CSA_sum_0_34_5, CSA_carry_0_34_5, CSA_sum_0_34_6, CSA_carry_0_34_6, CSA_sum_0_34_7, CSA_carry_0_34_7, CSA_sum_0_34_8, CSA_carry_0_34_8, CSA_sum_0_35_0, CSA_carry_0_35_0, CSA_sum_0_35_1, CSA_carry_0_35_1, CSA_sum_0_35_2, CSA_carry_0_35_2, CSA_sum_0_35_3, CSA_carry_0_35_3, CSA_sum_0_35_4, CSA_carry_0_35_4, CSA_sum_0_35_5, CSA_carry_0_35_5, CSA_sum_0_35_6, CSA_carry_0_35_6, CSA_sum_0_35_7, CSA_carry_0_35_7, CSA_sum_0_35_8, CSA_carry_0_35_8, CSA_sum_0_36_0, CSA_carry_0_36_0, CSA_sum_0_36_1, CSA_carry_0_36_1, CSA_sum_0_36_2, CSA_carry_0_36_2, CSA_sum_0_36_3, CSA_carry_0_36_3, CSA_sum_0_36_4, CSA_carry_0_36_4, CSA_sum_0_36_5, CSA_carry_0_36_5, CSA_sum_0_36_6, CSA_carry_0_36_6, CSA_sum_0_36_7, CSA_carry_0_36_7, CSA_sum_0_36_8, CSA_carry_0_36_8, CSA_sum_0_37_0, CSA_carry_0_37_0, CSA_sum_0_37_1, CSA_carry_0_37_1, CSA_sum_0_37_2, CSA_carry_0_37_2, CSA_sum_0_37_3, CSA_carry_0_37_3, CSA_sum_0_37_4, CSA_carry_0_37_4, CSA_sum_0_37_5, CSA_carry_0_37_5, CSA_sum_0_37_6, CSA_carry_0_37_6, CSA_sum_0_37_7, CSA_carry_0_37_7, CSA_sum_0_38_0, CSA_carry_0_38_0, CSA_sum_0_38_1, CSA_carry_0_38_1, CSA_sum_0_38_2, CSA_carry_0_38_2, CSA_sum_0_38_3, CSA_carry_0_38_3, CSA_sum_0_38_4, CSA_carry_0_38_4, CSA_sum_0_38_5, CSA_carry_0_38_5, CSA_sum_0_38_6, CSA_carry_0_38_6, CSA_sum_0_38_7, CSA_carry_0_38_7, CSA_sum_0_39_0, CSA_carry_0_39_0, CSA_sum_0_39_1, CSA_carry_0_39_1, CSA_sum_0_39_2, CSA_carry_0_39_2, CSA_sum_0_39_3, CSA_carry_0_39_3, CSA_sum_0_39_4, CSA_carry_0_39_4, CSA_sum_0_39_5, CSA_carry_0_39_5, CSA_sum_0_39_6, CSA_carry_0_39_6, CSA_sum_0_39_7, CSA_carry_0_39_7, CSA_sum_0_40_0, CSA_carry_0_40_0, CSA_sum_0_40_1, CSA_carry_0_40_1, CSA_sum_0_40_2, CSA_carry_0_40_2, CSA_sum_0_40_3, CSA_carry_0_40_3, CSA_sum_0_40_4, CSA_carry_0_40_4, CSA_sum_0_40_5, CSA_carry_0_40_5, CSA_sum_0_40_6, CSA_carry_0_40_6, CSA_sum_0_41_0, CSA_carry_0_41_0, CSA_sum_0_41_1, CSA_carry_0_41_1, CSA_sum_0_41_2, CSA_carry_0_41_2, CSA_sum_0_41_3, CSA_carry_0_41_3, CSA_sum_0_41_4, CSA_carry_0_41_4, CSA_sum_0_41_5, CSA_carry_0_41_5, CSA_sum_0_41_6, CSA_carry_0_41_6, CSA_sum_0_42_0, CSA_carry_0_42_0, CSA_sum_0_42_1, CSA_carry_0_42_1, CSA_sum_0_42_2, CSA_carry_0_42_2, CSA_sum_0_42_3, CSA_carry_0_42_3, CSA_sum_0_42_4, CSA_carry_0_42_4, CSA_sum_0_42_5, CSA_carry_0_42_5, CSA_sum_0_42_6, CSA_carry_0_42_6, CSA_sum_0_43_0, CSA_carry_0_43_0, CSA_sum_0_43_1, CSA_carry_0_43_1, CSA_sum_0_43_2, CSA_carry_0_43_2, CSA_sum_0_43_3, CSA_carry_0_43_3, CSA_sum_0_43_4, CSA_carry_0_43_4, CSA_sum_0_43_5, CSA_carry_0_43_5, CSA_sum_0_44_0, CSA_carry_0_44_0, CSA_sum_0_44_1, CSA_carry_0_44_1, CSA_sum_0_44_2, CSA_carry_0_44_2, CSA_sum_0_44_3, CSA_carry_0_44_3, CSA_sum_0_44_4, CSA_carry_0_44_4, CSA_sum_0_44_5, CSA_carry_0_44_5, CSA_sum_0_45_0, CSA_carry_0_45_0, CSA_sum_0_45_1, CSA_carry_0_45_1, CSA_sum_0_45_2, CSA_carry_0_45_2, CSA_sum_0_45_3, CSA_carry_0_45_3, CSA_sum_0_45_4, CSA_carry_0_45_4, CSA_sum_0_45_5, CSA_carry_0_45_5, CSA_sum_0_46_0, CSA_carry_0_46_0, CSA_sum_0_46_1, CSA_carry_0_46_1, CSA_sum_0_46_2, CSA_carry_0_46_2, CSA_sum_0_46_3, CSA_carry_0_46_3, CSA_sum_0_46_4, CSA_carry_0_46_4, CSA_sum_0_47_0, CSA_carry_0_47_0, CSA_sum_0_47_1, CSA_carry_0_47_1, CSA_sum_0_47_2, CSA_carry_0_47_2, CSA_sum_0_47_3, CSA_carry_0_47_3, CSA_sum_0_47_4, CSA_carry_0_47_4, CSA_sum_0_48_0, CSA_carry_0_48_0, CSA_sum_0_48_1, CSA_carry_0_48_1, CSA_sum_0_48_2, CSA_carry_0_48_2, CSA_sum_0_48_3, CSA_carry_0_48_3, CSA_sum_0_48_4, CSA_carry_0_48_4, CSA_sum_0_49_0, CSA_carry_0_49_0, CSA_sum_0_49_1, CSA_carry_0_49_1, CSA_sum_0_49_2, CSA_carry_0_49_2, CSA_sum_0_49_3, CSA_carry_0_49_3, CSA_sum_0_50_0, CSA_carry_0_50_0, CSA_sum_0_50_1, CSA_carry_0_50_1, CSA_sum_0_50_2, CSA_carry_0_50_2, CSA_sum_0_50_3, CSA_carry_0_50_3, CSA_sum_0_51_0, CSA_carry_0_51_0, CSA_sum_0_51_1, CSA_carry_0_51_1, CSA_sum_0_51_2, CSA_carry_0_51_2, CSA_sum_0_51_3, CSA_carry_0_51_3, CSA_sum_0_52_0, CSA_carry_0_52_0, CSA_sum_0_52_1, CSA_carry_0_52_1, CSA_sum_0_52_2, CSA_carry_0_52_2, CSA_sum_0_53_0, CSA_carry_0_53_0, CSA_sum_0_53_1, CSA_carry_0_53_1, CSA_sum_0_53_2, CSA_carry_0_53_2, CSA_sum_0_54_0, CSA_carry_0_54_0, CSA_sum_0_54_1, CSA_carry_0_54_1, CSA_sum_0_54_2, CSA_carry_0_54_2, CSA_sum_0_55_0, CSA_carry_0_55_0, CSA_sum_0_55_1, CSA_carry_0_55_1, CSA_sum_0_56_0, CSA_carry_0_56_0, CSA_sum_0_56_1, CSA_carry_0_56_1, CSA_sum_0_57_0, CSA_carry_0_57_0, CSA_sum_0_57_1, CSA_carry_0_57_1, CSA_sum_0_58_0, CSA_carry_0_58_0, CSA_sum_0_59_0, CSA_carry_0_59_0, CSA_sum_0_60_0, CSA_carry_0_60_0 : std_logic;
--signals for iteration 1
signal CSA_sum_1_3_0, CSA_carry_1_3_0, CSA_sum_1_4_0, CSA_carry_1_4_0, CSA_sum_1_5_0, CSA_carry_1_5_0, CSA_sum_1_6_0, CSA_carry_1_6_0, CSA_sum_1_7_0, CSA_carry_1_7_0, CSA_sum_1_7_1, CSA_carry_1_7_1, CSA_sum_1_8_0, CSA_carry_1_8_0, CSA_sum_1_9_0, CSA_carry_1_9_0, CSA_sum_1_9_1, CSA_carry_1_9_1, CSA_sum_1_10_0, CSA_carry_1_10_0, CSA_sum_1_10_1, CSA_carry_1_10_1, CSA_sum_1_11_0, CSA_carry_1_11_0, CSA_sum_1_11_1, CSA_carry_1_11_1, CSA_sum_1_12_0, CSA_carry_1_12_0, CSA_sum_1_12_1, CSA_carry_1_12_1, CSA_sum_1_12_2, CSA_carry_1_12_2, CSA_sum_1_13_0, CSA_carry_1_13_0, CSA_sum_1_13_1, CSA_carry_1_13_1, CSA_sum_1_13_2, CSA_carry_1_13_2, CSA_sum_1_14_0, CSA_carry_1_14_0, CSA_sum_1_14_1, CSA_carry_1_14_1, CSA_sum_1_14_2, CSA_carry_1_14_2, CSA_sum_1_15_0, CSA_carry_1_15_0, CSA_sum_1_15_1, CSA_carry_1_15_1, CSA_sum_1_15_2, CSA_carry_1_15_2, CSA_sum_1_16_0, CSA_carry_1_16_0, CSA_sum_1_16_1, CSA_carry_1_16_1, CSA_sum_1_16_2, CSA_carry_1_16_2, CSA_sum_1_16_3, CSA_carry_1_16_3, CSA_sum_1_17_0, CSA_carry_1_17_0, CSA_sum_1_17_1, CSA_carry_1_17_1, CSA_sum_1_17_2, CSA_carry_1_17_2, CSA_sum_1_18_0, CSA_carry_1_18_0, CSA_sum_1_18_1, CSA_carry_1_18_1, CSA_sum_1_18_2, CSA_carry_1_18_2, CSA_sum_1_18_3, CSA_carry_1_18_3, CSA_sum_1_19_0, CSA_carry_1_19_0, CSA_sum_1_19_1, CSA_carry_1_19_1, CSA_sum_1_19_2, CSA_carry_1_19_2, CSA_sum_1_19_3, CSA_carry_1_19_3, CSA_sum_1_20_0, CSA_carry_1_20_0, CSA_sum_1_20_1, CSA_carry_1_20_1, CSA_sum_1_20_2, CSA_carry_1_20_2, CSA_sum_1_20_3, CSA_carry_1_20_3, CSA_sum_1_21_0, CSA_carry_1_21_0, CSA_sum_1_21_1, CSA_carry_1_21_1, CSA_sum_1_21_2, CSA_carry_1_21_2, CSA_sum_1_21_3, CSA_carry_1_21_3, CSA_sum_1_21_4, CSA_carry_1_21_4, CSA_sum_1_22_0, CSA_carry_1_22_0, CSA_sum_1_22_1, CSA_carry_1_22_1, CSA_sum_1_22_2, CSA_carry_1_22_2, CSA_sum_1_22_3, CSA_carry_1_22_3, CSA_sum_1_22_4, CSA_carry_1_22_4, CSA_sum_1_23_0, CSA_carry_1_23_0, CSA_sum_1_23_1, CSA_carry_1_23_1, CSA_sum_1_23_2, CSA_carry_1_23_2, CSA_sum_1_23_3, CSA_carry_1_23_3, CSA_sum_1_23_4, CSA_carry_1_23_4, CSA_sum_1_24_0, CSA_carry_1_24_0, CSA_sum_1_24_1, CSA_carry_1_24_1, CSA_sum_1_24_2, CSA_carry_1_24_2, CSA_sum_1_24_3, CSA_carry_1_24_3, CSA_sum_1_24_4, CSA_carry_1_24_4, CSA_sum_1_25_0, CSA_carry_1_25_0, CSA_sum_1_25_1, CSA_carry_1_25_1, CSA_sum_1_25_2, CSA_carry_1_25_2, CSA_sum_1_25_3, CSA_carry_1_25_3, CSA_sum_1_25_4, CSA_carry_1_25_4, CSA_sum_1_25_5, CSA_carry_1_25_5, CSA_sum_1_26_0, CSA_carry_1_26_0, CSA_sum_1_26_1, CSA_carry_1_26_1, CSA_sum_1_26_2, CSA_carry_1_26_2, CSA_sum_1_26_3, CSA_carry_1_26_3, CSA_sum_1_26_4, CSA_carry_1_26_4, CSA_sum_1_27_0, CSA_carry_1_27_0, CSA_sum_1_27_1, CSA_carry_1_27_1, CSA_sum_1_27_2, CSA_carry_1_27_2, CSA_sum_1_27_3, CSA_carry_1_27_3, CSA_sum_1_27_4, CSA_carry_1_27_4, CSA_sum_1_27_5, CSA_carry_1_27_5, CSA_sum_1_28_0, CSA_carry_1_28_0, CSA_sum_1_28_1, CSA_carry_1_28_1, CSA_sum_1_28_2, CSA_carry_1_28_2, CSA_sum_1_28_3, CSA_carry_1_28_3, CSA_sum_1_28_4, CSA_carry_1_28_4, CSA_sum_1_28_5, CSA_carry_1_28_5, CSA_sum_1_29_0, CSA_carry_1_29_0, CSA_sum_1_29_1, CSA_carry_1_29_1, CSA_sum_1_29_2, CSA_carry_1_29_2, CSA_sum_1_29_3, CSA_carry_1_29_3, CSA_sum_1_29_4, CSA_carry_1_29_4, CSA_sum_1_29_5, CSA_carry_1_29_5, CSA_sum_1_30_0, CSA_carry_1_30_0, CSA_sum_1_30_1, CSA_carry_1_30_1, CSA_sum_1_30_2, CSA_carry_1_30_2, CSA_sum_1_30_3, CSA_carry_1_30_3, CSA_sum_1_30_4, CSA_carry_1_30_4, CSA_sum_1_30_5, CSA_carry_1_30_5, CSA_sum_1_30_6, CSA_carry_1_30_6, CSA_sum_1_31_0, CSA_carry_1_31_0, CSA_sum_1_31_1, CSA_carry_1_31_1, CSA_sum_1_31_2, CSA_carry_1_31_2, CSA_sum_1_31_3, CSA_carry_1_31_3, CSA_sum_1_31_4, CSA_carry_1_31_4, CSA_sum_1_31_5, CSA_carry_1_31_5, CSA_sum_1_31_6, CSA_carry_1_31_6, CSA_sum_1_32_0, CSA_carry_1_32_0, CSA_sum_1_32_1, CSA_carry_1_32_1, CSA_sum_1_32_2, CSA_carry_1_32_2, CSA_sum_1_32_3, CSA_carry_1_32_3, CSA_sum_1_32_4, CSA_carry_1_32_4, CSA_sum_1_32_5, CSA_carry_1_32_5, CSA_sum_1_32_6, CSA_carry_1_32_6, CSA_sum_1_33_0, CSA_carry_1_33_0, CSA_sum_1_33_1, CSA_carry_1_33_1, CSA_sum_1_33_2, CSA_carry_1_33_2, CSA_sum_1_33_3, CSA_carry_1_33_3, CSA_sum_1_33_4, CSA_carry_1_33_4, CSA_sum_1_33_5, CSA_carry_1_33_5, CSA_sum_1_34_0, CSA_carry_1_34_0, CSA_sum_1_34_1, CSA_carry_1_34_1, CSA_sum_1_34_2, CSA_carry_1_34_2, CSA_sum_1_34_3, CSA_carry_1_34_3, CSA_sum_1_34_4, CSA_carry_1_34_4, CSA_sum_1_34_5, CSA_carry_1_34_5, CSA_sum_1_34_6, CSA_carry_1_34_6, CSA_sum_1_35_0, CSA_carry_1_35_0, CSA_sum_1_35_1, CSA_carry_1_35_1, CSA_sum_1_35_2, CSA_carry_1_35_2, CSA_sum_1_35_3, CSA_carry_1_35_3, CSA_sum_1_35_4, CSA_carry_1_35_4, CSA_sum_1_35_5, CSA_carry_1_35_5, CSA_sum_1_36_0, CSA_carry_1_36_0, CSA_sum_1_36_1, CSA_carry_1_36_1, CSA_sum_1_36_2, CSA_carry_1_36_2, CSA_sum_1_36_3, CSA_carry_1_36_3, CSA_sum_1_36_4, CSA_carry_1_36_4, CSA_sum_1_36_5, CSA_carry_1_36_5, CSA_sum_1_37_0, CSA_carry_1_37_0, CSA_sum_1_37_1, CSA_carry_1_37_1, CSA_sum_1_37_2, CSA_carry_1_37_2, CSA_sum_1_37_3, CSA_carry_1_37_3, CSA_sum_1_37_4, CSA_carry_1_37_4, CSA_sum_1_37_5, CSA_carry_1_37_5, CSA_sum_1_38_0, CSA_carry_1_38_0, CSA_sum_1_38_1, CSA_carry_1_38_1, CSA_sum_1_38_2, CSA_carry_1_38_2, CSA_sum_1_38_3, CSA_carry_1_38_3, CSA_sum_1_38_4, CSA_carry_1_38_4, CSA_sum_1_39_0, CSA_carry_1_39_0, CSA_sum_1_39_1, CSA_carry_1_39_1, CSA_sum_1_39_2, CSA_carry_1_39_2, CSA_sum_1_39_3, CSA_carry_1_39_3, CSA_sum_1_39_4, CSA_carry_1_39_4, CSA_sum_1_40_0, CSA_carry_1_40_0, CSA_sum_1_40_1, CSA_carry_1_40_1, CSA_sum_1_40_2, CSA_carry_1_40_2, CSA_sum_1_40_3, CSA_carry_1_40_3, CSA_sum_1_40_4, CSA_carry_1_40_4, CSA_sum_1_41_0, CSA_carry_1_41_0, CSA_sum_1_41_1, CSA_carry_1_41_1, CSA_sum_1_41_2, CSA_carry_1_41_2, CSA_sum_1_41_3, CSA_carry_1_41_3, CSA_sum_1_41_4, CSA_carry_1_41_4, CSA_sum_1_42_0, CSA_carry_1_42_0, CSA_sum_1_42_1, CSA_carry_1_42_1, CSA_sum_1_42_2, CSA_carry_1_42_2, CSA_sum_1_42_3, CSA_carry_1_42_3, CSA_sum_1_43_0, CSA_carry_1_43_0, CSA_sum_1_43_1, CSA_carry_1_43_1, CSA_sum_1_43_2, CSA_carry_1_43_2, CSA_sum_1_43_3, CSA_carry_1_43_3, CSA_sum_1_43_4, CSA_carry_1_43_4, CSA_sum_1_44_0, CSA_carry_1_44_0, CSA_sum_1_44_1, CSA_carry_1_44_1, CSA_sum_1_44_2, CSA_carry_1_44_2, CSA_sum_1_44_3, CSA_carry_1_44_3, CSA_sum_1_45_0, CSA_carry_1_45_0, CSA_sum_1_45_1, CSA_carry_1_45_1, CSA_sum_1_45_2, CSA_carry_1_45_2, CSA_sum_1_45_3, CSA_carry_1_45_3, CSA_sum_1_46_0, CSA_carry_1_46_0, CSA_sum_1_46_1, CSA_carry_1_46_1, CSA_sum_1_46_2, CSA_carry_1_46_2, CSA_sum_1_46_3, CSA_carry_1_46_3, CSA_sum_1_47_0, CSA_carry_1_47_0, CSA_sum_1_47_1, CSA_carry_1_47_1, CSA_sum_1_47_2, CSA_carry_1_47_2, CSA_sum_1_48_0, CSA_carry_1_48_0, CSA_sum_1_48_1, CSA_carry_1_48_1, CSA_sum_1_48_2, CSA_carry_1_48_2, CSA_sum_1_49_0, CSA_carry_1_49_0, CSA_sum_1_49_1, CSA_carry_1_49_1, CSA_sum_1_49_2, CSA_carry_1_49_2, CSA_sum_1_50_0, CSA_carry_1_50_0, CSA_sum_1_50_1, CSA_carry_1_50_1, CSA_sum_1_50_2, CSA_carry_1_50_2, CSA_sum_1_51_0, CSA_carry_1_51_0, CSA_sum_1_51_1, CSA_carry_1_51_1, CSA_sum_1_52_0, CSA_carry_1_52_0, CSA_sum_1_52_1, CSA_carry_1_52_1, CSA_sum_1_52_2, CSA_carry_1_52_2, CSA_sum_1_53_0, CSA_carry_1_53_0, CSA_sum_1_53_1, CSA_carry_1_53_1, CSA_sum_1_54_0, CSA_carry_1_54_0, CSA_sum_1_54_1, CSA_carry_1_54_1, CSA_sum_1_55_0, CSA_carry_1_55_0, CSA_sum_1_55_1, CSA_carry_1_55_1, CSA_sum_1_56_0, CSA_carry_1_56_0, CSA_sum_1_57_0, CSA_carry_1_57_0, CSA_sum_1_58_0, CSA_carry_1_58_0, CSA_sum_1_59_0, CSA_carry_1_59_0, CSA_sum_1_61_0, CSA_carry_1_61_0 : std_logic;
--signals for iteration 2
signal CSA_sum_2_4_0, CSA_carry_2_4_0, CSA_sum_2_6_0, CSA_carry_2_6_0, CSA_sum_2_7_0, CSA_carry_2_7_0, CSA_sum_2_8_0, CSA_carry_2_8_0, CSA_sum_2_9_0, CSA_carry_2_9_0, CSA_sum_2_10_0, CSA_carry_2_10_0, CSA_sum_2_10_1, CSA_carry_2_10_1, CSA_sum_2_11_0, CSA_carry_2_11_0, CSA_sum_2_12_0, CSA_carry_2_12_0, CSA_sum_2_13_0, CSA_carry_2_13_0, CSA_sum_2_13_1, CSA_carry_2_13_1, CSA_sum_2_14_0, CSA_carry_2_14_0, CSA_sum_2_14_1, CSA_carry_2_14_1, CSA_sum_2_15_0, CSA_carry_2_15_0, CSA_sum_2_15_1, CSA_carry_2_15_1, CSA_sum_2_16_0, CSA_carry_2_16_0, CSA_sum_2_16_1, CSA_carry_2_16_1, CSA_sum_2_17_0, CSA_carry_2_17_0, CSA_sum_2_17_1, CSA_carry_2_17_1, CSA_sum_2_17_2, CSA_carry_2_17_2, CSA_sum_2_18_0, CSA_carry_2_18_0, CSA_sum_2_18_1, CSA_carry_2_18_1, CSA_sum_2_19_0, CSA_carry_2_19_0, CSA_sum_2_19_1, CSA_carry_2_19_1, CSA_sum_2_19_2, CSA_carry_2_19_2, CSA_sum_2_20_0, CSA_carry_2_20_0, CSA_sum_2_20_1, CSA_carry_2_20_1, CSA_sum_2_20_2, CSA_carry_2_20_2, CSA_sum_2_21_0, CSA_carry_2_21_0, CSA_sum_2_21_1, CSA_carry_2_21_1, CSA_sum_2_21_2, CSA_carry_2_21_2, CSA_sum_2_22_0, CSA_carry_2_22_0, CSA_sum_2_22_1, CSA_carry_2_22_1, CSA_sum_2_22_2, CSA_carry_2_22_2, CSA_sum_2_23_0, CSA_carry_2_23_0, CSA_sum_2_23_1, CSA_carry_2_23_1, CSA_sum_2_23_2, CSA_carry_2_23_2, CSA_sum_2_24_0, CSA_carry_2_24_0, CSA_sum_2_24_1, CSA_carry_2_24_1, CSA_sum_2_24_2, CSA_carry_2_24_2, CSA_sum_2_24_3, CSA_carry_2_24_3, CSA_sum_2_25_0, CSA_carry_2_25_0, CSA_sum_2_25_1, CSA_carry_2_25_1, CSA_sum_2_25_2, CSA_carry_2_25_2, CSA_sum_2_26_0, CSA_carry_2_26_0, CSA_sum_2_26_1, CSA_carry_2_26_1, CSA_sum_2_26_2, CSA_carry_2_26_2, CSA_sum_2_26_3, CSA_carry_2_26_3, CSA_sum_2_27_0, CSA_carry_2_27_0, CSA_sum_2_27_1, CSA_carry_2_27_1, CSA_sum_2_27_2, CSA_carry_2_27_2, CSA_sum_2_27_3, CSA_carry_2_27_3, CSA_sum_2_28_0, CSA_carry_2_28_0, CSA_sum_2_28_1, CSA_carry_2_28_1, CSA_sum_2_28_2, CSA_carry_2_28_2, CSA_sum_2_28_3, CSA_carry_2_28_3, CSA_sum_2_29_0, CSA_carry_2_29_0, CSA_sum_2_29_1, CSA_carry_2_29_1, CSA_sum_2_29_2, CSA_carry_2_29_2, CSA_sum_2_29_3, CSA_carry_2_29_3, CSA_sum_2_30_0, CSA_carry_2_30_0, CSA_sum_2_30_1, CSA_carry_2_30_1, CSA_sum_2_30_2, CSA_carry_2_30_2, CSA_sum_2_30_3, CSA_carry_2_30_3, CSA_sum_2_31_0, CSA_carry_2_31_0, CSA_sum_2_31_1, CSA_carry_2_31_1, CSA_sum_2_31_2, CSA_carry_2_31_2, CSA_sum_2_31_3, CSA_carry_2_31_3, CSA_sum_2_31_4, CSA_carry_2_31_4, CSA_sum_2_32_0, CSA_carry_2_32_0, CSA_sum_2_32_1, CSA_carry_2_32_1, CSA_sum_2_32_2, CSA_carry_2_32_2, CSA_sum_2_32_3, CSA_carry_2_32_3, CSA_sum_2_33_0, CSA_carry_2_33_0, CSA_sum_2_33_1, CSA_carry_2_33_1, CSA_sum_2_33_2, CSA_carry_2_33_2, CSA_sum_2_33_3, CSA_carry_2_33_3, CSA_sum_2_33_4, CSA_carry_2_33_4, CSA_sum_2_34_0, CSA_carry_2_34_0, CSA_sum_2_34_1, CSA_carry_2_34_1, CSA_sum_2_34_2, CSA_carry_2_34_2, CSA_sum_2_34_3, CSA_carry_2_34_3, CSA_sum_2_35_0, CSA_carry_2_35_0, CSA_sum_2_35_1, CSA_carry_2_35_1, CSA_sum_2_35_2, CSA_carry_2_35_2, CSA_sum_2_35_3, CSA_carry_2_35_3, CSA_sum_2_36_0, CSA_carry_2_36_0, CSA_sum_2_36_1, CSA_carry_2_36_1, CSA_sum_2_36_2, CSA_carry_2_36_2, CSA_sum_2_36_3, CSA_carry_2_36_3, CSA_sum_2_37_0, CSA_carry_2_37_0, CSA_sum_2_37_1, CSA_carry_2_37_1, CSA_sum_2_37_2, CSA_carry_2_37_2, CSA_sum_2_37_3, CSA_carry_2_37_3, CSA_sum_2_38_0, CSA_carry_2_38_0, CSA_sum_2_38_1, CSA_carry_2_38_1, CSA_sum_2_38_2, CSA_carry_2_38_2, CSA_sum_2_38_3, CSA_carry_2_38_3, CSA_sum_2_39_0, CSA_carry_2_39_0, CSA_sum_2_39_1, CSA_carry_2_39_1, CSA_sum_2_39_2, CSA_carry_2_39_2, CSA_sum_2_40_0, CSA_carry_2_40_0, CSA_sum_2_40_1, CSA_carry_2_40_1, CSA_sum_2_40_2, CSA_carry_2_40_2, CSA_sum_2_40_3, CSA_carry_2_40_3, CSA_sum_2_41_0, CSA_carry_2_41_0, CSA_sum_2_41_1, CSA_carry_2_41_1, CSA_sum_2_41_2, CSA_carry_2_41_2, CSA_sum_2_42_0, CSA_carry_2_42_0, CSA_sum_2_42_1, CSA_carry_2_42_1, CSA_sum_2_42_2, CSA_carry_2_42_2, CSA_sum_2_43_0, CSA_carry_2_43_0, CSA_sum_2_43_1, CSA_carry_2_43_1, CSA_sum_2_43_2, CSA_carry_2_43_2, CSA_sum_2_44_0, CSA_carry_2_44_0, CSA_sum_2_44_1, CSA_carry_2_44_1, CSA_sum_2_44_2, CSA_carry_2_44_2, CSA_sum_2_45_0, CSA_carry_2_45_0, CSA_sum_2_45_1, CSA_carry_2_45_1, CSA_sum_2_46_0, CSA_carry_2_46_0, CSA_sum_2_46_1, CSA_carry_2_46_1, CSA_sum_2_46_2, CSA_carry_2_46_2, CSA_sum_2_47_0, CSA_carry_2_47_0, CSA_sum_2_47_1, CSA_carry_2_47_1, CSA_sum_2_47_2, CSA_carry_2_47_2, CSA_sum_2_48_0, CSA_carry_2_48_0, CSA_sum_2_48_1, CSA_carry_2_48_1, CSA_sum_2_49_0, CSA_carry_2_49_0, CSA_sum_2_49_1, CSA_carry_2_49_1, CSA_sum_2_50_0, CSA_carry_2_50_0, CSA_sum_2_50_1, CSA_carry_2_50_1, CSA_sum_2_51_0, CSA_carry_2_51_0, CSA_sum_2_51_1, CSA_carry_2_51_1, CSA_sum_2_52_0, CSA_carry_2_52_0, CSA_sum_2_53_0, CSA_carry_2_53_0, CSA_sum_2_53_1, CSA_carry_2_53_1, CSA_sum_2_54_0, CSA_carry_2_54_0, CSA_sum_2_55_0, CSA_carry_2_55_0, CSA_sum_2_56_0, CSA_carry_2_56_0, CSA_sum_2_57_0, CSA_carry_2_57_0, CSA_sum_2_58_0, CSA_carry_2_58_0, CSA_sum_2_60_0, CSA_carry_2_60_0 : std_logic;
--signals for iteration 3
signal CSA_sum_3_5_0, CSA_carry_3_5_0, CSA_sum_3_8_0, CSA_carry_3_8_0, CSA_sum_3_9_0, CSA_carry_3_9_0, CSA_sum_3_10_0, CSA_carry_3_10_0, CSA_sum_3_11_0, CSA_carry_3_11_0, CSA_sum_3_12_0, CSA_carry_3_12_0, CSA_sum_3_13_0, CSA_carry_3_13_0, CSA_sum_3_14_0, CSA_carry_3_14_0, CSA_sum_3_15_0, CSA_carry_3_15_0, CSA_sum_3_15_1, CSA_carry_3_15_1, CSA_sum_3_16_0, CSA_carry_3_16_0, CSA_sum_3_17_0, CSA_carry_3_17_0, CSA_sum_3_18_0, CSA_carry_3_18_0, CSA_sum_3_18_1, CSA_carry_3_18_1, CSA_sum_3_19_0, CSA_carry_3_19_0, CSA_sum_3_19_1, CSA_carry_3_19_1, CSA_sum_3_20_0, CSA_carry_3_20_0, CSA_sum_3_20_1, CSA_carry_3_20_1, CSA_sum_3_21_0, CSA_carry_3_21_0, CSA_sum_3_21_1, CSA_carry_3_21_1, CSA_sum_3_22_0, CSA_carry_3_22_0, CSA_sum_3_22_1, CSA_carry_3_22_1, CSA_sum_3_23_0, CSA_carry_3_23_0, CSA_sum_3_23_1, CSA_carry_3_23_1, CSA_sum_3_24_0, CSA_carry_3_24_0, CSA_sum_3_24_1, CSA_carry_3_24_1, CSA_sum_3_25_0, CSA_carry_3_25_0, CSA_sum_3_25_1, CSA_carry_3_25_1, CSA_sum_3_25_2, CSA_carry_3_25_2, CSA_sum_3_26_0, CSA_carry_3_26_0, CSA_sum_3_26_1, CSA_carry_3_26_1, CSA_sum_3_27_0, CSA_carry_3_27_0, CSA_sum_3_27_1, CSA_carry_3_27_1, CSA_sum_3_28_0, CSA_carry_3_28_0, CSA_sum_3_28_1, CSA_carry_3_28_1, CSA_sum_3_28_2, CSA_carry_3_28_2, CSA_sum_3_29_0, CSA_carry_3_29_0, CSA_sum_3_29_1, CSA_carry_3_29_1, CSA_sum_3_29_2, CSA_carry_3_29_2, CSA_sum_3_30_0, CSA_carry_3_30_0, CSA_sum_3_30_1, CSA_carry_3_30_1, CSA_sum_3_30_2, CSA_carry_3_30_2, CSA_sum_3_31_0, CSA_carry_3_31_0, CSA_sum_3_31_1, CSA_carry_3_31_1, CSA_sum_3_31_2, CSA_carry_3_31_2, CSA_sum_3_32_0, CSA_carry_3_32_0, CSA_sum_3_32_1, CSA_carry_3_32_1, CSA_sum_3_32_2, CSA_carry_3_32_2, CSA_sum_3_33_0, CSA_carry_3_33_0, CSA_sum_3_33_1, CSA_carry_3_33_1, CSA_sum_3_33_2, CSA_carry_3_33_2, CSA_sum_3_34_0, CSA_carry_3_34_0, CSA_sum_3_34_1, CSA_carry_3_34_1, CSA_sum_3_34_2, CSA_carry_3_34_2, CSA_sum_3_35_0, CSA_carry_3_35_0, CSA_sum_3_35_1, CSA_carry_3_35_1, CSA_sum_3_35_2, CSA_carry_3_35_2, CSA_sum_3_36_0, CSA_carry_3_36_0, CSA_sum_3_36_1, CSA_carry_3_36_1, CSA_sum_3_37_0, CSA_carry_3_37_0, CSA_sum_3_37_1, CSA_carry_3_37_1, CSA_sum_3_37_2, CSA_carry_3_37_2, CSA_sum_3_38_0, CSA_carry_3_38_0, CSA_sum_3_38_1, CSA_carry_3_38_1, CSA_sum_3_38_2, CSA_carry_3_38_2, CSA_sum_3_39_0, CSA_carry_3_39_0, CSA_sum_3_39_1, CSA_carry_3_39_1, CSA_sum_3_39_2, CSA_carry_3_39_2, CSA_sum_3_40_0, CSA_carry_3_40_0, CSA_sum_3_40_1, CSA_carry_3_40_1, CSA_sum_3_41_0, CSA_carry_3_41_0, CSA_sum_3_41_1, CSA_carry_3_41_1, CSA_sum_3_42_0, CSA_carry_3_42_0, CSA_sum_3_42_1, CSA_carry_3_42_1, CSA_sum_3_43_0, CSA_carry_3_43_0, CSA_sum_3_43_1, CSA_carry_3_43_1, CSA_sum_3_44_0, CSA_carry_3_44_0, CSA_sum_3_44_1, CSA_carry_3_44_1, CSA_sum_3_45_0, CSA_carry_3_45_0, CSA_sum_3_45_1, CSA_carry_3_45_1, CSA_sum_3_46_0, CSA_carry_3_46_0, CSA_sum_3_47_0, CSA_carry_3_47_0, CSA_sum_3_47_1, CSA_carry_3_47_1, CSA_sum_3_48_0, CSA_carry_3_48_0, CSA_sum_3_48_1, CSA_carry_3_48_1, CSA_sum_3_49_0, CSA_carry_3_49_0, CSA_sum_3_49_1, CSA_carry_3_49_1, CSA_sum_3_50_0, CSA_carry_3_50_0, CSA_sum_3_51_0, CSA_carry_3_51_0, CSA_sum_3_52_0, CSA_carry_3_52_0, CSA_sum_3_53_0, CSA_carry_3_53_0, CSA_sum_3_54_0, CSA_carry_3_54_0, CSA_sum_3_55_0, CSA_carry_3_55_0, CSA_sum_3_56_0, CSA_carry_3_56_0, CSA_sum_3_58_0, CSA_carry_3_58_0, CSA_sum_3_59_0, CSA_carry_3_59_0 : std_logic;
--signals for iteration 4
signal CSA_sum_4_6_0, CSA_carry_4_6_0, CSA_sum_4_11_0, CSA_carry_4_11_0, CSA_sum_4_12_0, CSA_carry_4_12_0, CSA_sum_4_13_0, CSA_carry_4_13_0, CSA_sum_4_14_0, CSA_carry_4_14_0, CSA_sum_4_15_0, CSA_carry_4_15_0, CSA_sum_4_16_0, CSA_carry_4_16_0, CSA_sum_4_17_0, CSA_carry_4_17_0, CSA_sum_4_18_0, CSA_carry_4_18_0, CSA_sum_4_19_0, CSA_carry_4_19_0, CSA_sum_4_20_0, CSA_carry_4_20_0, CSA_sum_4_21_0, CSA_carry_4_21_0, CSA_sum_4_22_0, CSA_carry_4_22_0, CSA_sum_4_22_1, CSA_carry_4_22_1, CSA_sum_4_23_0, CSA_carry_4_23_0, CSA_sum_4_24_0, CSA_carry_4_24_0, CSA_sum_4_25_0, CSA_carry_4_25_0, CSA_sum_4_26_0, CSA_carry_4_26_0, CSA_sum_4_26_1, CSA_carry_4_26_1, CSA_sum_4_27_0, CSA_carry_4_27_0, CSA_sum_4_27_1, CSA_carry_4_27_1, CSA_sum_4_28_0, CSA_carry_4_28_0, CSA_sum_4_28_1, CSA_carry_4_28_1, CSA_sum_4_29_0, CSA_carry_4_29_0, CSA_sum_4_29_1, CSA_carry_4_29_1, CSA_sum_4_30_0, CSA_carry_4_30_0, CSA_sum_4_30_1, CSA_carry_4_30_1, CSA_sum_4_31_0, CSA_carry_4_31_0, CSA_sum_4_31_1, CSA_carry_4_31_1, CSA_sum_4_32_0, CSA_carry_4_32_0, CSA_sum_4_32_1, CSA_carry_4_32_1, CSA_sum_4_33_0, CSA_carry_4_33_0, CSA_sum_4_33_1, CSA_carry_4_33_1, CSA_sum_4_34_0, CSA_carry_4_34_0, CSA_sum_4_34_1, CSA_carry_4_34_1, CSA_sum_4_35_0, CSA_carry_4_35_0, CSA_sum_4_35_1, CSA_carry_4_35_1, CSA_sum_4_36_0, CSA_carry_4_36_0, CSA_sum_4_36_1, CSA_carry_4_36_1, CSA_sum_4_37_0, CSA_carry_4_37_0, CSA_sum_4_38_0, CSA_carry_4_38_0, CSA_sum_4_38_1, CSA_carry_4_38_1, CSA_sum_4_39_0, CSA_carry_4_39_0, CSA_sum_4_39_1, CSA_carry_4_39_1, CSA_sum_4_40_0, CSA_carry_4_40_0, CSA_sum_4_40_1, CSA_carry_4_40_1, CSA_sum_4_41_0, CSA_carry_4_41_0, CSA_sum_4_41_1, CSA_carry_4_41_1, CSA_sum_4_42_0, CSA_carry_4_42_0, CSA_sum_4_42_1, CSA_carry_4_42_1, CSA_sum_4_43_0, CSA_carry_4_43_0, CSA_sum_4_44_0, CSA_carry_4_44_0, CSA_sum_4_45_0, CSA_carry_4_45_0, CSA_sum_4_46_0, CSA_carry_4_46_0, CSA_sum_4_47_0, CSA_carry_4_47_0, CSA_sum_4_48_0, CSA_carry_4_48_0, CSA_sum_4_49_0, CSA_carry_4_49_0, CSA_sum_4_50_0, CSA_carry_4_50_0, CSA_sum_4_51_0, CSA_carry_4_51_0, CSA_sum_4_52_0, CSA_carry_4_52_0, CSA_sum_4_54_0, CSA_carry_4_54_0, CSA_sum_4_55_0, CSA_carry_4_55_0, CSA_sum_4_56_0, CSA_carry_4_56_0, CSA_sum_4_57_0, CSA_carry_4_57_0 : std_logic;
--signals for iteration 5
signal CSA_sum_5_7_0, CSA_carry_5_7_0, CSA_sum_5_16_0, CSA_carry_5_16_0, CSA_sum_5_17_0, CSA_carry_5_17_0, CSA_sum_5_18_0, CSA_carry_5_18_0, CSA_sum_5_19_0, CSA_carry_5_19_0, CSA_sum_5_20_0, CSA_carry_5_20_0, CSA_sum_5_21_0, CSA_carry_5_21_0, CSA_sum_5_22_0, CSA_carry_5_22_0, CSA_sum_5_23_0, CSA_carry_5_23_0, CSA_sum_5_24_0, CSA_carry_5_24_0, CSA_sum_5_25_0, CSA_carry_5_25_0, CSA_sum_5_26_0, CSA_carry_5_26_0, CSA_sum_5_27_0, CSA_carry_5_27_0, CSA_sum_5_28_0, CSA_carry_5_28_0, CSA_sum_5_29_0, CSA_carry_5_29_0, CSA_sum_5_30_0, CSA_carry_5_30_0, CSA_sum_5_31_0, CSA_carry_5_31_0, CSA_sum_5_32_0, CSA_carry_5_32_0, CSA_sum_5_32_1, CSA_carry_5_32_1, CSA_sum_5_33_0, CSA_carry_5_33_0, CSA_sum_5_34_0, CSA_carry_5_34_0, CSA_sum_5_35_0, CSA_carry_5_35_0, CSA_sum_5_36_0, CSA_carry_5_36_0, CSA_sum_5_37_0, CSA_carry_5_37_0, CSA_sum_5_38_0, CSA_carry_5_38_0, CSA_sum_5_39_0, CSA_carry_5_39_0, CSA_sum_5_40_0, CSA_carry_5_40_0, CSA_sum_5_41_0, CSA_carry_5_41_0, CSA_sum_5_42_0, CSA_carry_5_42_0, CSA_sum_5_43_0, CSA_carry_5_43_0, CSA_sum_5_44_0, CSA_carry_5_44_0, CSA_sum_5_45_0, CSA_carry_5_45_0, CSA_sum_5_46_0, CSA_carry_5_46_0, CSA_sum_5_48_0, CSA_carry_5_48_0, CSA_sum_5_49_0, CSA_carry_5_49_0, CSA_sum_5_50_0, CSA_carry_5_50_0, CSA_sum_5_51_0, CSA_carry_5_51_0, CSA_sum_5_52_0, CSA_carry_5_52_0, CSA_sum_5_53_0, CSA_carry_5_53_0 : std_logic;
--signals for iteration 6
signal CSA_sum_6_8_0, CSA_carry_6_8_0, CSA_sum_6_23_0, CSA_carry_6_23_0, CSA_sum_6_24_0, CSA_carry_6_24_0, CSA_sum_6_25_0, CSA_carry_6_25_0, CSA_sum_6_26_0, CSA_carry_6_26_0, CSA_sum_6_27_0, CSA_carry_6_27_0, CSA_sum_6_28_0, CSA_carry_6_28_0, CSA_sum_6_29_0, CSA_carry_6_29_0, CSA_sum_6_30_0, CSA_carry_6_30_0, CSA_sum_6_31_0, CSA_carry_6_31_0, CSA_sum_6_32_0, CSA_carry_6_32_0, CSA_sum_6_33_0, CSA_carry_6_33_0, CSA_sum_6_34_0, CSA_carry_6_34_0, CSA_sum_6_35_0, CSA_carry_6_35_0, CSA_sum_6_36_0, CSA_carry_6_36_0, CSA_sum_6_37_0, CSA_carry_6_37_0, CSA_sum_6_39_0, CSA_carry_6_39_0, CSA_sum_6_40_0, CSA_carry_6_40_0, CSA_sum_6_41_0, CSA_carry_6_41_0, CSA_sum_6_42_0, CSA_carry_6_42_0, CSA_sum_6_43_0, CSA_carry_6_43_0, CSA_sum_6_44_0, CSA_carry_6_44_0, CSA_sum_6_45_0, CSA_carry_6_45_0, CSA_sum_6_46_0, CSA_carry_6_46_0, CSA_sum_6_47_0, CSA_carry_6_47_0 : std_logic;
--signals for iteration 7
signal CSA_sum_7_9_0, CSA_carry_7_9_0, CSA_sum_7_33_0, CSA_carry_7_33_0, CSA_sum_7_34_0, CSA_carry_7_34_0, CSA_sum_7_35_0, CSA_carry_7_35_0, CSA_sum_7_36_0, CSA_carry_7_36_0, CSA_sum_7_37_0, CSA_carry_7_37_0, CSA_sum_7_38_0, CSA_carry_7_38_0 : std_logic;
--signals for iteration 8
signal CSA_sum_8_10_0, CSA_carry_8_10_0 : std_logic;
--signals for iteration 9
signal CSA_sum_9_11_0, CSA_carry_9_11_0 : std_logic;
--signals for iteration 10
signal CSA_sum_10_12_0, CSA_carry_10_12_0 : std_logic;
--signals for iteration 11
signal CSA_sum_11_13_0, CSA_carry_11_13_0 : std_logic;
--signals for iteration 12
signal CSA_sum_12_14_0, CSA_carry_12_14_0 : std_logic;
--signals for iteration 13
signal CSA_sum_13_15_0, CSA_carry_13_15_0 : std_logic;
--signals for iteration 14
signal CSA_sum_14_16_0, CSA_carry_14_16_0 : std_logic;
--signals for iteration 15
signal CSA_sum_15_17_0, CSA_carry_15_17_0 : std_logic;
--signals for iteration 16
signal CSA_sum_16_18_0, CSA_carry_16_18_0 : std_logic;
--signals for iteration 17
signal CSA_sum_17_19_0, CSA_carry_17_19_0 : std_logic;
--signals for iteration 18
signal CSA_sum_18_20_0, CSA_carry_18_20_0 : std_logic;
--signals for iteration 19
signal CSA_sum_19_21_0, CSA_carry_19_21_0 : std_logic;
--signals for iteration 20
signal CSA_sum_20_22_0, CSA_carry_20_22_0 : std_logic;
--signals for iteration 21
signal CSA_sum_21_23_0, CSA_carry_21_23_0 : std_logic;
--signals for iteration 22
signal CSA_sum_22_24_0, CSA_carry_22_24_0 : std_logic;
--signals for iteration 23
signal CSA_sum_23_25_0, CSA_carry_23_25_0 : std_logic;
--signals for iteration 24
signal CSA_sum_24_26_0, CSA_carry_24_26_0 : std_logic;
--signals for iteration 25
signal CSA_sum_25_27_0, CSA_carry_25_27_0 : std_logic;
--signals for iteration 26
signal CSA_sum_26_28_0, CSA_carry_26_28_0 : std_logic;
--signals for iteration 27
signal CSA_sum_27_29_0, CSA_carry_27_29_0 : std_logic;
--signals for iteration 28
signal CSA_sum_28_30_0, CSA_carry_28_30_0 : std_logic;
--signals for iteration 29
signal CSA_sum_29_31_0, CSA_carry_29_31_0 : std_logic;
--signals for iteration 30
signal CSA_sum_30_32_0, CSA_carry_30_32_0 : std_logic;

signal b_and_a : std_logic_vector(1023 downto 0);
begin

gen3: for X in 31 downto 0 generate
gen4X: for Y in 31 downto 0 generate
b_and_a(X + 32*Y) <= in1(X) AND in2(Y);
end generate;
end generate;
FA_lbl_0_2_0: FA port map(in1 => b_and_a(2), in2 => b_and_a(33), c_in => b_and_a(64), sum => CSA_sum_0_2_0, c_out => CSA_carry_0_2_0);
FA_lbl_0_3_0: FA port map(in1 => b_and_a(3), in2 => b_and_a(34), c_in => b_and_a(65), sum => CSA_sum_0_3_0, c_out => CSA_carry_0_3_0);
FA_lbl_0_4_0: FA port map(in1 => b_and_a(4), in2 => b_and_a(35), c_in => b_and_a(66), sum => CSA_sum_0_4_0, c_out => CSA_carry_0_4_0);
FA_lbl_0_5_0: FA port map(in1 => b_and_a(5), in2 => b_and_a(36), c_in => b_and_a(67), sum => CSA_sum_0_5_0, c_out => CSA_carry_0_5_0);
FA_lbl_0_5_1: FA port map(in1 => b_and_a(98), in2 => b_and_a(129), c_in => b_and_a(160), sum => CSA_sum_0_5_1, c_out => CSA_carry_0_5_1);
FA_lbl_0_6_0: FA port map(in1 => b_and_a(6), in2 => b_and_a(37), c_in => b_and_a(68), sum => CSA_sum_0_6_0, c_out => CSA_carry_0_6_0);
FA_lbl_0_6_1: FA port map(in1 => b_and_a(99), in2 => b_and_a(130), c_in => b_and_a(161), sum => CSA_sum_0_6_1, c_out => CSA_carry_0_6_1);
FA_lbl_0_7_0: FA port map(in1 => b_and_a(7), in2 => b_and_a(38), c_in => b_and_a(69), sum => CSA_sum_0_7_0, c_out => CSA_carry_0_7_0);
FA_lbl_0_7_1: FA port map(in1 => b_and_a(100), in2 => b_and_a(131), c_in => b_and_a(162), sum => CSA_sum_0_7_1, c_out => CSA_carry_0_7_1);
FA_lbl_0_8_0: FA port map(in1 => b_and_a(8), in2 => b_and_a(39), c_in => b_and_a(70), sum => CSA_sum_0_8_0, c_out => CSA_carry_0_8_0);
FA_lbl_0_8_1: FA port map(in1 => b_and_a(101), in2 => b_and_a(132), c_in => b_and_a(163), sum => CSA_sum_0_8_1, c_out => CSA_carry_0_8_1);
FA_lbl_0_8_2: FA port map(in1 => b_and_a(194), in2 => b_and_a(225), c_in => b_and_a(256), sum => CSA_sum_0_8_2, c_out => CSA_carry_0_8_2);
FA_lbl_0_9_0: FA port map(in1 => b_and_a(9), in2 => b_and_a(40), c_in => b_and_a(71), sum => CSA_sum_0_9_0, c_out => CSA_carry_0_9_0);
FA_lbl_0_9_1: FA port map(in1 => b_and_a(102), in2 => b_and_a(133), c_in => b_and_a(164), sum => CSA_sum_0_9_1, c_out => CSA_carry_0_9_1);
FA_lbl_0_9_2: FA port map(in1 => b_and_a(195), in2 => b_and_a(226), c_in => b_and_a(257), sum => CSA_sum_0_9_2, c_out => CSA_carry_0_9_2);
FA_lbl_0_10_0: FA port map(in1 => b_and_a(10), in2 => b_and_a(41), c_in => b_and_a(72), sum => CSA_sum_0_10_0, c_out => CSA_carry_0_10_0);
FA_lbl_0_10_1: FA port map(in1 => b_and_a(103), in2 => b_and_a(134), c_in => b_and_a(165), sum => CSA_sum_0_10_1, c_out => CSA_carry_0_10_1);
FA_lbl_0_10_2: FA port map(in1 => b_and_a(196), in2 => b_and_a(227), c_in => b_and_a(258), sum => CSA_sum_0_10_2, c_out => CSA_carry_0_10_2);
FA_lbl_0_11_0: FA port map(in1 => b_and_a(11), in2 => b_and_a(42), c_in => b_and_a(73), sum => CSA_sum_0_11_0, c_out => CSA_carry_0_11_0);
FA_lbl_0_11_1: FA port map(in1 => b_and_a(104), in2 => b_and_a(135), c_in => b_and_a(166), sum => CSA_sum_0_11_1, c_out => CSA_carry_0_11_1);
FA_lbl_0_11_2: FA port map(in1 => b_and_a(197), in2 => b_and_a(228), c_in => b_and_a(259), sum => CSA_sum_0_11_2, c_out => CSA_carry_0_11_2);
FA_lbl_0_11_3: FA port map(in1 => b_and_a(290), in2 => b_and_a(321), c_in => b_and_a(352), sum => CSA_sum_0_11_3, c_out => CSA_carry_0_11_3);
FA_lbl_0_12_0: FA port map(in1 => b_and_a(12), in2 => b_and_a(43), c_in => b_and_a(74), sum => CSA_sum_0_12_0, c_out => CSA_carry_0_12_0);
FA_lbl_0_12_1: FA port map(in1 => b_and_a(105), in2 => b_and_a(136), c_in => b_and_a(167), sum => CSA_sum_0_12_1, c_out => CSA_carry_0_12_1);
FA_lbl_0_12_2: FA port map(in1 => b_and_a(198), in2 => b_and_a(229), c_in => b_and_a(260), sum => CSA_sum_0_12_2, c_out => CSA_carry_0_12_2);
FA_lbl_0_12_3: FA port map(in1 => b_and_a(291), in2 => b_and_a(322), c_in => b_and_a(353), sum => CSA_sum_0_12_3, c_out => CSA_carry_0_12_3);
FA_lbl_0_13_0: FA port map(in1 => b_and_a(13), in2 => b_and_a(44), c_in => b_and_a(75), sum => CSA_sum_0_13_0, c_out => CSA_carry_0_13_0);
FA_lbl_0_13_1: FA port map(in1 => b_and_a(106), in2 => b_and_a(137), c_in => b_and_a(168), sum => CSA_sum_0_13_1, c_out => CSA_carry_0_13_1);
FA_lbl_0_13_2: FA port map(in1 => b_and_a(199), in2 => b_and_a(230), c_in => b_and_a(261), sum => CSA_sum_0_13_2, c_out => CSA_carry_0_13_2);
FA_lbl_0_13_3: FA port map(in1 => b_and_a(292), in2 => b_and_a(323), c_in => b_and_a(354), sum => CSA_sum_0_13_3, c_out => CSA_carry_0_13_3);
FA_lbl_0_14_0: FA port map(in1 => b_and_a(14), in2 => b_and_a(45), c_in => b_and_a(76), sum => CSA_sum_0_14_0, c_out => CSA_carry_0_14_0);
FA_lbl_0_14_1: FA port map(in1 => b_and_a(107), in2 => b_and_a(138), c_in => b_and_a(169), sum => CSA_sum_0_14_1, c_out => CSA_carry_0_14_1);
FA_lbl_0_14_2: FA port map(in1 => b_and_a(200), in2 => b_and_a(231), c_in => b_and_a(262), sum => CSA_sum_0_14_2, c_out => CSA_carry_0_14_2);
FA_lbl_0_14_3: FA port map(in1 => b_and_a(293), in2 => b_and_a(324), c_in => b_and_a(355), sum => CSA_sum_0_14_3, c_out => CSA_carry_0_14_3);
FA_lbl_0_14_4: FA port map(in1 => b_and_a(386), in2 => b_and_a(417), c_in => b_and_a(448), sum => CSA_sum_0_14_4, c_out => CSA_carry_0_14_4);
FA_lbl_0_15_0: FA port map(in1 => b_and_a(15), in2 => b_and_a(46), c_in => b_and_a(77), sum => CSA_sum_0_15_0, c_out => CSA_carry_0_15_0);
FA_lbl_0_15_1: FA port map(in1 => b_and_a(108), in2 => b_and_a(139), c_in => b_and_a(170), sum => CSA_sum_0_15_1, c_out => CSA_carry_0_15_1);
FA_lbl_0_15_2: FA port map(in1 => b_and_a(201), in2 => b_and_a(232), c_in => b_and_a(263), sum => CSA_sum_0_15_2, c_out => CSA_carry_0_15_2);
FA_lbl_0_15_3: FA port map(in1 => b_and_a(294), in2 => b_and_a(325), c_in => b_and_a(356), sum => CSA_sum_0_15_3, c_out => CSA_carry_0_15_3);
FA_lbl_0_15_4: FA port map(in1 => b_and_a(387), in2 => b_and_a(418), c_in => b_and_a(449), sum => CSA_sum_0_15_4, c_out => CSA_carry_0_15_4);
FA_lbl_0_16_0: FA port map(in1 => b_and_a(16), in2 => b_and_a(47), c_in => b_and_a(78), sum => CSA_sum_0_16_0, c_out => CSA_carry_0_16_0);
FA_lbl_0_16_1: FA port map(in1 => b_and_a(109), in2 => b_and_a(140), c_in => b_and_a(171), sum => CSA_sum_0_16_1, c_out => CSA_carry_0_16_1);
FA_lbl_0_16_2: FA port map(in1 => b_and_a(202), in2 => b_and_a(233), c_in => b_and_a(264), sum => CSA_sum_0_16_2, c_out => CSA_carry_0_16_2);
FA_lbl_0_16_3: FA port map(in1 => b_and_a(295), in2 => b_and_a(326), c_in => b_and_a(357), sum => CSA_sum_0_16_3, c_out => CSA_carry_0_16_3);
FA_lbl_0_16_4: FA port map(in1 => b_and_a(388), in2 => b_and_a(419), c_in => b_and_a(450), sum => CSA_sum_0_16_4, c_out => CSA_carry_0_16_4);
FA_lbl_0_17_0: FA port map(in1 => b_and_a(17), in2 => b_and_a(48), c_in => b_and_a(79), sum => CSA_sum_0_17_0, c_out => CSA_carry_0_17_0);
FA_lbl_0_17_1: FA port map(in1 => b_and_a(110), in2 => b_and_a(141), c_in => b_and_a(172), sum => CSA_sum_0_17_1, c_out => CSA_carry_0_17_1);
FA_lbl_0_17_2: FA port map(in1 => b_and_a(203), in2 => b_and_a(234), c_in => b_and_a(265), sum => CSA_sum_0_17_2, c_out => CSA_carry_0_17_2);
FA_lbl_0_17_3: FA port map(in1 => b_and_a(296), in2 => b_and_a(327), c_in => b_and_a(358), sum => CSA_sum_0_17_3, c_out => CSA_carry_0_17_3);
FA_lbl_0_17_4: FA port map(in1 => b_and_a(389), in2 => b_and_a(420), c_in => b_and_a(451), sum => CSA_sum_0_17_4, c_out => CSA_carry_0_17_4);
FA_lbl_0_17_5: FA port map(in1 => b_and_a(482), in2 => b_and_a(513), c_in => b_and_a(544), sum => CSA_sum_0_17_5, c_out => CSA_carry_0_17_5);
FA_lbl_0_18_0: FA port map(in1 => b_and_a(18), in2 => b_and_a(49), c_in => b_and_a(80), sum => CSA_sum_0_18_0, c_out => CSA_carry_0_18_0);
FA_lbl_0_18_1: FA port map(in1 => b_and_a(111), in2 => b_and_a(142), c_in => b_and_a(173), sum => CSA_sum_0_18_1, c_out => CSA_carry_0_18_1);
FA_lbl_0_18_2: FA port map(in1 => b_and_a(204), in2 => b_and_a(235), c_in => b_and_a(266), sum => CSA_sum_0_18_2, c_out => CSA_carry_0_18_2);
FA_lbl_0_18_3: FA port map(in1 => b_and_a(297), in2 => b_and_a(328), c_in => b_and_a(359), sum => CSA_sum_0_18_3, c_out => CSA_carry_0_18_3);
FA_lbl_0_18_4: FA port map(in1 => b_and_a(390), in2 => b_and_a(421), c_in => b_and_a(452), sum => CSA_sum_0_18_4, c_out => CSA_carry_0_18_4);
FA_lbl_0_18_5: FA port map(in1 => b_and_a(483), in2 => b_and_a(514), c_in => b_and_a(545), sum => CSA_sum_0_18_5, c_out => CSA_carry_0_18_5);
FA_lbl_0_19_0: FA port map(in1 => b_and_a(19), in2 => b_and_a(50), c_in => b_and_a(81), sum => CSA_sum_0_19_0, c_out => CSA_carry_0_19_0);
FA_lbl_0_19_1: FA port map(in1 => b_and_a(112), in2 => b_and_a(143), c_in => b_and_a(174), sum => CSA_sum_0_19_1, c_out => CSA_carry_0_19_1);
FA_lbl_0_19_2: FA port map(in1 => b_and_a(205), in2 => b_and_a(236), c_in => b_and_a(267), sum => CSA_sum_0_19_2, c_out => CSA_carry_0_19_2);
FA_lbl_0_19_3: FA port map(in1 => b_and_a(298), in2 => b_and_a(329), c_in => b_and_a(360), sum => CSA_sum_0_19_3, c_out => CSA_carry_0_19_3);
FA_lbl_0_19_4: FA port map(in1 => b_and_a(391), in2 => b_and_a(422), c_in => b_and_a(453), sum => CSA_sum_0_19_4, c_out => CSA_carry_0_19_4);
FA_lbl_0_19_5: FA port map(in1 => b_and_a(484), in2 => b_and_a(515), c_in => b_and_a(546), sum => CSA_sum_0_19_5, c_out => CSA_carry_0_19_5);
FA_lbl_0_20_0: FA port map(in1 => b_and_a(20), in2 => b_and_a(51), c_in => b_and_a(82), sum => CSA_sum_0_20_0, c_out => CSA_carry_0_20_0);
FA_lbl_0_20_1: FA port map(in1 => b_and_a(113), in2 => b_and_a(144), c_in => b_and_a(175), sum => CSA_sum_0_20_1, c_out => CSA_carry_0_20_1);
FA_lbl_0_20_2: FA port map(in1 => b_and_a(206), in2 => b_and_a(237), c_in => b_and_a(268), sum => CSA_sum_0_20_2, c_out => CSA_carry_0_20_2);
FA_lbl_0_20_3: FA port map(in1 => b_and_a(299), in2 => b_and_a(330), c_in => b_and_a(361), sum => CSA_sum_0_20_3, c_out => CSA_carry_0_20_3);
FA_lbl_0_20_4: FA port map(in1 => b_and_a(392), in2 => b_and_a(423), c_in => b_and_a(454), sum => CSA_sum_0_20_4, c_out => CSA_carry_0_20_4);
FA_lbl_0_20_5: FA port map(in1 => b_and_a(485), in2 => b_and_a(516), c_in => b_and_a(547), sum => CSA_sum_0_20_5, c_out => CSA_carry_0_20_5);
FA_lbl_0_20_6: FA port map(in1 => b_and_a(578), in2 => b_and_a(609), c_in => b_and_a(640), sum => CSA_sum_0_20_6, c_out => CSA_carry_0_20_6);
FA_lbl_0_21_0: FA port map(in1 => b_and_a(21), in2 => b_and_a(52), c_in => b_and_a(83), sum => CSA_sum_0_21_0, c_out => CSA_carry_0_21_0);
FA_lbl_0_21_1: FA port map(in1 => b_and_a(114), in2 => b_and_a(145), c_in => b_and_a(176), sum => CSA_sum_0_21_1, c_out => CSA_carry_0_21_1);
FA_lbl_0_21_2: FA port map(in1 => b_and_a(207), in2 => b_and_a(238), c_in => b_and_a(269), sum => CSA_sum_0_21_2, c_out => CSA_carry_0_21_2);
FA_lbl_0_21_3: FA port map(in1 => b_and_a(300), in2 => b_and_a(331), c_in => b_and_a(362), sum => CSA_sum_0_21_3, c_out => CSA_carry_0_21_3);
FA_lbl_0_21_4: FA port map(in1 => b_and_a(393), in2 => b_and_a(424), c_in => b_and_a(455), sum => CSA_sum_0_21_4, c_out => CSA_carry_0_21_4);
FA_lbl_0_21_5: FA port map(in1 => b_and_a(486), in2 => b_and_a(517), c_in => b_and_a(548), sum => CSA_sum_0_21_5, c_out => CSA_carry_0_21_5);
FA_lbl_0_21_6: FA port map(in1 => b_and_a(579), in2 => b_and_a(610), c_in => b_and_a(641), sum => CSA_sum_0_21_6, c_out => CSA_carry_0_21_6);
FA_lbl_0_22_0: FA port map(in1 => b_and_a(22), in2 => b_and_a(53), c_in => b_and_a(84), sum => CSA_sum_0_22_0, c_out => CSA_carry_0_22_0);
FA_lbl_0_22_1: FA port map(in1 => b_and_a(115), in2 => b_and_a(146), c_in => b_and_a(177), sum => CSA_sum_0_22_1, c_out => CSA_carry_0_22_1);
FA_lbl_0_22_2: FA port map(in1 => b_and_a(208), in2 => b_and_a(239), c_in => b_and_a(270), sum => CSA_sum_0_22_2, c_out => CSA_carry_0_22_2);
FA_lbl_0_22_3: FA port map(in1 => b_and_a(301), in2 => b_and_a(332), c_in => b_and_a(363), sum => CSA_sum_0_22_3, c_out => CSA_carry_0_22_3);
FA_lbl_0_22_4: FA port map(in1 => b_and_a(394), in2 => b_and_a(425), c_in => b_and_a(456), sum => CSA_sum_0_22_4, c_out => CSA_carry_0_22_4);
FA_lbl_0_22_5: FA port map(in1 => b_and_a(487), in2 => b_and_a(518), c_in => b_and_a(549), sum => CSA_sum_0_22_5, c_out => CSA_carry_0_22_5);
FA_lbl_0_22_6: FA port map(in1 => b_and_a(580), in2 => b_and_a(611), c_in => b_and_a(642), sum => CSA_sum_0_22_6, c_out => CSA_carry_0_22_6);
FA_lbl_0_23_0: FA port map(in1 => b_and_a(23), in2 => b_and_a(54), c_in => b_and_a(85), sum => CSA_sum_0_23_0, c_out => CSA_carry_0_23_0);
FA_lbl_0_23_1: FA port map(in1 => b_and_a(116), in2 => b_and_a(147), c_in => b_and_a(178), sum => CSA_sum_0_23_1, c_out => CSA_carry_0_23_1);
FA_lbl_0_23_2: FA port map(in1 => b_and_a(209), in2 => b_and_a(240), c_in => b_and_a(271), sum => CSA_sum_0_23_2, c_out => CSA_carry_0_23_2);
FA_lbl_0_23_3: FA port map(in1 => b_and_a(302), in2 => b_and_a(333), c_in => b_and_a(364), sum => CSA_sum_0_23_3, c_out => CSA_carry_0_23_3);
FA_lbl_0_23_4: FA port map(in1 => b_and_a(395), in2 => b_and_a(426), c_in => b_and_a(457), sum => CSA_sum_0_23_4, c_out => CSA_carry_0_23_4);
FA_lbl_0_23_5: FA port map(in1 => b_and_a(488), in2 => b_and_a(519), c_in => b_and_a(550), sum => CSA_sum_0_23_5, c_out => CSA_carry_0_23_5);
FA_lbl_0_23_6: FA port map(in1 => b_and_a(581), in2 => b_and_a(612), c_in => b_and_a(643), sum => CSA_sum_0_23_6, c_out => CSA_carry_0_23_6);
FA_lbl_0_23_7: FA port map(in1 => b_and_a(674), in2 => b_and_a(705), c_in => b_and_a(736), sum => CSA_sum_0_23_7, c_out => CSA_carry_0_23_7);
FA_lbl_0_24_0: FA port map(in1 => b_and_a(24), in2 => b_and_a(55), c_in => b_and_a(86), sum => CSA_sum_0_24_0, c_out => CSA_carry_0_24_0);
FA_lbl_0_24_1: FA port map(in1 => b_and_a(117), in2 => b_and_a(148), c_in => b_and_a(179), sum => CSA_sum_0_24_1, c_out => CSA_carry_0_24_1);
FA_lbl_0_24_2: FA port map(in1 => b_and_a(210), in2 => b_and_a(241), c_in => b_and_a(272), sum => CSA_sum_0_24_2, c_out => CSA_carry_0_24_2);
FA_lbl_0_24_3: FA port map(in1 => b_and_a(303), in2 => b_and_a(334), c_in => b_and_a(365), sum => CSA_sum_0_24_3, c_out => CSA_carry_0_24_3);
FA_lbl_0_24_4: FA port map(in1 => b_and_a(396), in2 => b_and_a(427), c_in => b_and_a(458), sum => CSA_sum_0_24_4, c_out => CSA_carry_0_24_4);
FA_lbl_0_24_5: FA port map(in1 => b_and_a(489), in2 => b_and_a(520), c_in => b_and_a(551), sum => CSA_sum_0_24_5, c_out => CSA_carry_0_24_5);
FA_lbl_0_24_6: FA port map(in1 => b_and_a(582), in2 => b_and_a(613), c_in => b_and_a(644), sum => CSA_sum_0_24_6, c_out => CSA_carry_0_24_6);
FA_lbl_0_24_7: FA port map(in1 => b_and_a(675), in2 => b_and_a(706), c_in => b_and_a(737), sum => CSA_sum_0_24_7, c_out => CSA_carry_0_24_7);
FA_lbl_0_25_0: FA port map(in1 => b_and_a(25), in2 => b_and_a(56), c_in => b_and_a(87), sum => CSA_sum_0_25_0, c_out => CSA_carry_0_25_0);
FA_lbl_0_25_1: FA port map(in1 => b_and_a(118), in2 => b_and_a(149), c_in => b_and_a(180), sum => CSA_sum_0_25_1, c_out => CSA_carry_0_25_1);
FA_lbl_0_25_2: FA port map(in1 => b_and_a(211), in2 => b_and_a(242), c_in => b_and_a(273), sum => CSA_sum_0_25_2, c_out => CSA_carry_0_25_2);
FA_lbl_0_25_3: FA port map(in1 => b_and_a(304), in2 => b_and_a(335), c_in => b_and_a(366), sum => CSA_sum_0_25_3, c_out => CSA_carry_0_25_3);
FA_lbl_0_25_4: FA port map(in1 => b_and_a(397), in2 => b_and_a(428), c_in => b_and_a(459), sum => CSA_sum_0_25_4, c_out => CSA_carry_0_25_4);
FA_lbl_0_25_5: FA port map(in1 => b_and_a(490), in2 => b_and_a(521), c_in => b_and_a(552), sum => CSA_sum_0_25_5, c_out => CSA_carry_0_25_5);
FA_lbl_0_25_6: FA port map(in1 => b_and_a(583), in2 => b_and_a(614), c_in => b_and_a(645), sum => CSA_sum_0_25_6, c_out => CSA_carry_0_25_6);
FA_lbl_0_25_7: FA port map(in1 => b_and_a(676), in2 => b_and_a(707), c_in => b_and_a(738), sum => CSA_sum_0_25_7, c_out => CSA_carry_0_25_7);
FA_lbl_0_26_0: FA port map(in1 => b_and_a(26), in2 => b_and_a(57), c_in => b_and_a(88), sum => CSA_sum_0_26_0, c_out => CSA_carry_0_26_0);
FA_lbl_0_26_1: FA port map(in1 => b_and_a(119), in2 => b_and_a(150), c_in => b_and_a(181), sum => CSA_sum_0_26_1, c_out => CSA_carry_0_26_1);
FA_lbl_0_26_2: FA port map(in1 => b_and_a(212), in2 => b_and_a(243), c_in => b_and_a(274), sum => CSA_sum_0_26_2, c_out => CSA_carry_0_26_2);
FA_lbl_0_26_3: FA port map(in1 => b_and_a(305), in2 => b_and_a(336), c_in => b_and_a(367), sum => CSA_sum_0_26_3, c_out => CSA_carry_0_26_3);
FA_lbl_0_26_4: FA port map(in1 => b_and_a(398), in2 => b_and_a(429), c_in => b_and_a(460), sum => CSA_sum_0_26_4, c_out => CSA_carry_0_26_4);
FA_lbl_0_26_5: FA port map(in1 => b_and_a(491), in2 => b_and_a(522), c_in => b_and_a(553), sum => CSA_sum_0_26_5, c_out => CSA_carry_0_26_5);
FA_lbl_0_26_6: FA port map(in1 => b_and_a(584), in2 => b_and_a(615), c_in => b_and_a(646), sum => CSA_sum_0_26_6, c_out => CSA_carry_0_26_6);
FA_lbl_0_26_7: FA port map(in1 => b_and_a(677), in2 => b_and_a(708), c_in => b_and_a(739), sum => CSA_sum_0_26_7, c_out => CSA_carry_0_26_7);
FA_lbl_0_26_8: FA port map(in1 => b_and_a(770), in2 => b_and_a(801), c_in => b_and_a(832), sum => CSA_sum_0_26_8, c_out => CSA_carry_0_26_8);
FA_lbl_0_27_0: FA port map(in1 => b_and_a(27), in2 => b_and_a(58), c_in => b_and_a(89), sum => CSA_sum_0_27_0, c_out => CSA_carry_0_27_0);
FA_lbl_0_27_1: FA port map(in1 => b_and_a(120), in2 => b_and_a(151), c_in => b_and_a(182), sum => CSA_sum_0_27_1, c_out => CSA_carry_0_27_1);
FA_lbl_0_27_2: FA port map(in1 => b_and_a(213), in2 => b_and_a(244), c_in => b_and_a(275), sum => CSA_sum_0_27_2, c_out => CSA_carry_0_27_2);
FA_lbl_0_27_3: FA port map(in1 => b_and_a(306), in2 => b_and_a(337), c_in => b_and_a(368), sum => CSA_sum_0_27_3, c_out => CSA_carry_0_27_3);
FA_lbl_0_27_4: FA port map(in1 => b_and_a(399), in2 => b_and_a(430), c_in => b_and_a(461), sum => CSA_sum_0_27_4, c_out => CSA_carry_0_27_4);
FA_lbl_0_27_5: FA port map(in1 => b_and_a(492), in2 => b_and_a(523), c_in => b_and_a(554), sum => CSA_sum_0_27_5, c_out => CSA_carry_0_27_5);
FA_lbl_0_27_6: FA port map(in1 => b_and_a(585), in2 => b_and_a(616), c_in => b_and_a(647), sum => CSA_sum_0_27_6, c_out => CSA_carry_0_27_6);
FA_lbl_0_27_7: FA port map(in1 => b_and_a(678), in2 => b_and_a(709), c_in => b_and_a(740), sum => CSA_sum_0_27_7, c_out => CSA_carry_0_27_7);
FA_lbl_0_27_8: FA port map(in1 => b_and_a(771), in2 => b_and_a(802), c_in => b_and_a(833), sum => CSA_sum_0_27_8, c_out => CSA_carry_0_27_8);
FA_lbl_0_28_0: FA port map(in1 => b_and_a(28), in2 => b_and_a(59), c_in => b_and_a(90), sum => CSA_sum_0_28_0, c_out => CSA_carry_0_28_0);
FA_lbl_0_28_1: FA port map(in1 => b_and_a(121), in2 => b_and_a(152), c_in => b_and_a(183), sum => CSA_sum_0_28_1, c_out => CSA_carry_0_28_1);
FA_lbl_0_28_2: FA port map(in1 => b_and_a(214), in2 => b_and_a(245), c_in => b_and_a(276), sum => CSA_sum_0_28_2, c_out => CSA_carry_0_28_2);
FA_lbl_0_28_3: FA port map(in1 => b_and_a(307), in2 => b_and_a(338), c_in => b_and_a(369), sum => CSA_sum_0_28_3, c_out => CSA_carry_0_28_3);
FA_lbl_0_28_4: FA port map(in1 => b_and_a(400), in2 => b_and_a(431), c_in => b_and_a(462), sum => CSA_sum_0_28_4, c_out => CSA_carry_0_28_4);
FA_lbl_0_28_5: FA port map(in1 => b_and_a(493), in2 => b_and_a(524), c_in => b_and_a(555), sum => CSA_sum_0_28_5, c_out => CSA_carry_0_28_5);
FA_lbl_0_28_6: FA port map(in1 => b_and_a(586), in2 => b_and_a(617), c_in => b_and_a(648), sum => CSA_sum_0_28_6, c_out => CSA_carry_0_28_6);
FA_lbl_0_28_7: FA port map(in1 => b_and_a(679), in2 => b_and_a(710), c_in => b_and_a(741), sum => CSA_sum_0_28_7, c_out => CSA_carry_0_28_7);
FA_lbl_0_28_8: FA port map(in1 => b_and_a(772), in2 => b_and_a(803), c_in => b_and_a(834), sum => CSA_sum_0_28_8, c_out => CSA_carry_0_28_8);
FA_lbl_0_29_0: FA port map(in1 => b_and_a(29), in2 => b_and_a(60), c_in => b_and_a(91), sum => CSA_sum_0_29_0, c_out => CSA_carry_0_29_0);
FA_lbl_0_29_1: FA port map(in1 => b_and_a(122), in2 => b_and_a(153), c_in => b_and_a(184), sum => CSA_sum_0_29_1, c_out => CSA_carry_0_29_1);
FA_lbl_0_29_2: FA port map(in1 => b_and_a(215), in2 => b_and_a(246), c_in => b_and_a(277), sum => CSA_sum_0_29_2, c_out => CSA_carry_0_29_2);
FA_lbl_0_29_3: FA port map(in1 => b_and_a(308), in2 => b_and_a(339), c_in => b_and_a(370), sum => CSA_sum_0_29_3, c_out => CSA_carry_0_29_3);
FA_lbl_0_29_4: FA port map(in1 => b_and_a(401), in2 => b_and_a(432), c_in => b_and_a(463), sum => CSA_sum_0_29_4, c_out => CSA_carry_0_29_4);
FA_lbl_0_29_5: FA port map(in1 => b_and_a(494), in2 => b_and_a(525), c_in => b_and_a(556), sum => CSA_sum_0_29_5, c_out => CSA_carry_0_29_5);
FA_lbl_0_29_6: FA port map(in1 => b_and_a(587), in2 => b_and_a(618), c_in => b_and_a(649), sum => CSA_sum_0_29_6, c_out => CSA_carry_0_29_6);
FA_lbl_0_29_7: FA port map(in1 => b_and_a(680), in2 => b_and_a(711), c_in => b_and_a(742), sum => CSA_sum_0_29_7, c_out => CSA_carry_0_29_7);
FA_lbl_0_29_8: FA port map(in1 => b_and_a(773), in2 => b_and_a(804), c_in => b_and_a(835), sum => CSA_sum_0_29_8, c_out => CSA_carry_0_29_8);
FA_lbl_0_29_9: FA port map(in1 => b_and_a(866), in2 => b_and_a(897), c_in => b_and_a(928), sum => CSA_sum_0_29_9, c_out => CSA_carry_0_29_9);
FA_lbl_0_30_0: FA port map(in1 => b_and_a(30), in2 => b_and_a(61), c_in => b_and_a(92), sum => CSA_sum_0_30_0, c_out => CSA_carry_0_30_0);
FA_lbl_0_30_1: FA port map(in1 => b_and_a(123), in2 => b_and_a(154), c_in => b_and_a(185), sum => CSA_sum_0_30_1, c_out => CSA_carry_0_30_1);
FA_lbl_0_30_2: FA port map(in1 => b_and_a(216), in2 => b_and_a(247), c_in => b_and_a(278), sum => CSA_sum_0_30_2, c_out => CSA_carry_0_30_2);
FA_lbl_0_30_3: FA port map(in1 => b_and_a(309), in2 => b_and_a(340), c_in => b_and_a(371), sum => CSA_sum_0_30_3, c_out => CSA_carry_0_30_3);
FA_lbl_0_30_4: FA port map(in1 => b_and_a(402), in2 => b_and_a(433), c_in => b_and_a(464), sum => CSA_sum_0_30_4, c_out => CSA_carry_0_30_4);
FA_lbl_0_30_5: FA port map(in1 => b_and_a(495), in2 => b_and_a(526), c_in => b_and_a(557), sum => CSA_sum_0_30_5, c_out => CSA_carry_0_30_5);
FA_lbl_0_30_6: FA port map(in1 => b_and_a(588), in2 => b_and_a(619), c_in => b_and_a(650), sum => CSA_sum_0_30_6, c_out => CSA_carry_0_30_6);
FA_lbl_0_30_7: FA port map(in1 => b_and_a(681), in2 => b_and_a(712), c_in => b_and_a(743), sum => CSA_sum_0_30_7, c_out => CSA_carry_0_30_7);
FA_lbl_0_30_8: FA port map(in1 => b_and_a(774), in2 => b_and_a(805), c_in => b_and_a(836), sum => CSA_sum_0_30_8, c_out => CSA_carry_0_30_8);
FA_lbl_0_30_9: FA port map(in1 => b_and_a(867), in2 => b_and_a(898), c_in => b_and_a(929), sum => CSA_sum_0_30_9, c_out => CSA_carry_0_30_9);
FA_lbl_0_31_0: FA port map(in1 => b_and_a(31), in2 => b_and_a(62), c_in => b_and_a(93), sum => CSA_sum_0_31_0, c_out => CSA_carry_0_31_0);
FA_lbl_0_31_1: FA port map(in1 => b_and_a(124), in2 => b_and_a(155), c_in => b_and_a(186), sum => CSA_sum_0_31_1, c_out => CSA_carry_0_31_1);
FA_lbl_0_31_2: FA port map(in1 => b_and_a(217), in2 => b_and_a(248), c_in => b_and_a(279), sum => CSA_sum_0_31_2, c_out => CSA_carry_0_31_2);
FA_lbl_0_31_3: FA port map(in1 => b_and_a(310), in2 => b_and_a(341), c_in => b_and_a(372), sum => CSA_sum_0_31_3, c_out => CSA_carry_0_31_3);
FA_lbl_0_31_4: FA port map(in1 => b_and_a(403), in2 => b_and_a(434), c_in => b_and_a(465), sum => CSA_sum_0_31_4, c_out => CSA_carry_0_31_4);
FA_lbl_0_31_5: FA port map(in1 => b_and_a(496), in2 => b_and_a(527), c_in => b_and_a(558), sum => CSA_sum_0_31_5, c_out => CSA_carry_0_31_5);
FA_lbl_0_31_6: FA port map(in1 => b_and_a(589), in2 => b_and_a(620), c_in => b_and_a(651), sum => CSA_sum_0_31_6, c_out => CSA_carry_0_31_6);
FA_lbl_0_31_7: FA port map(in1 => b_and_a(682), in2 => b_and_a(713), c_in => b_and_a(744), sum => CSA_sum_0_31_7, c_out => CSA_carry_0_31_7);
FA_lbl_0_31_8: FA port map(in1 => b_and_a(775), in2 => b_and_a(806), c_in => b_and_a(837), sum => CSA_sum_0_31_8, c_out => CSA_carry_0_31_8);
FA_lbl_0_31_9: FA port map(in1 => b_and_a(868), in2 => b_and_a(899), c_in => b_and_a(930), sum => CSA_sum_0_31_9, c_out => CSA_carry_0_31_9);
FA_lbl_0_32_0: FA port map(in1 => b_and_a(63), in2 => b_and_a(94), c_in => b_and_a(125), sum => CSA_sum_0_32_0, c_out => CSA_carry_0_32_0);
FA_lbl_0_32_1: FA port map(in1 => b_and_a(156), in2 => b_and_a(187), c_in => b_and_a(218), sum => CSA_sum_0_32_1, c_out => CSA_carry_0_32_1);
FA_lbl_0_32_2: FA port map(in1 => b_and_a(249), in2 => b_and_a(280), c_in => b_and_a(311), sum => CSA_sum_0_32_2, c_out => CSA_carry_0_32_2);
FA_lbl_0_32_3: FA port map(in1 => b_and_a(342), in2 => b_and_a(373), c_in => b_and_a(404), sum => CSA_sum_0_32_3, c_out => CSA_carry_0_32_3);
FA_lbl_0_32_4: FA port map(in1 => b_and_a(435), in2 => b_and_a(466), c_in => b_and_a(497), sum => CSA_sum_0_32_4, c_out => CSA_carry_0_32_4);
FA_lbl_0_32_5: FA port map(in1 => b_and_a(528), in2 => b_and_a(559), c_in => b_and_a(590), sum => CSA_sum_0_32_5, c_out => CSA_carry_0_32_5);
FA_lbl_0_32_6: FA port map(in1 => b_and_a(621), in2 => b_and_a(652), c_in => b_and_a(683), sum => CSA_sum_0_32_6, c_out => CSA_carry_0_32_6);
FA_lbl_0_32_7: FA port map(in1 => b_and_a(714), in2 => b_and_a(745), c_in => b_and_a(776), sum => CSA_sum_0_32_7, c_out => CSA_carry_0_32_7);
FA_lbl_0_32_8: FA port map(in1 => b_and_a(807), in2 => b_and_a(838), c_in => b_and_a(869), sum => CSA_sum_0_32_8, c_out => CSA_carry_0_32_8);
FA_lbl_0_32_9: FA port map(in1 => b_and_a(900), in2 => b_and_a(931), c_in => b_and_a(962), sum => CSA_sum_0_32_9, c_out => CSA_carry_0_32_9);
FA_lbl_0_33_0: FA port map(in1 => b_and_a(95), in2 => b_and_a(126), c_in => b_and_a(157), sum => CSA_sum_0_33_0, c_out => CSA_carry_0_33_0);
FA_lbl_0_33_1: FA port map(in1 => b_and_a(188), in2 => b_and_a(219), c_in => b_and_a(250), sum => CSA_sum_0_33_1, c_out => CSA_carry_0_33_1);
FA_lbl_0_33_2: FA port map(in1 => b_and_a(281), in2 => b_and_a(312), c_in => b_and_a(343), sum => CSA_sum_0_33_2, c_out => CSA_carry_0_33_2);
FA_lbl_0_33_3: FA port map(in1 => b_and_a(374), in2 => b_and_a(405), c_in => b_and_a(436), sum => CSA_sum_0_33_3, c_out => CSA_carry_0_33_3);
FA_lbl_0_33_4: FA port map(in1 => b_and_a(467), in2 => b_and_a(498), c_in => b_and_a(529), sum => CSA_sum_0_33_4, c_out => CSA_carry_0_33_4);
FA_lbl_0_33_5: FA port map(in1 => b_and_a(560), in2 => b_and_a(591), c_in => b_and_a(622), sum => CSA_sum_0_33_5, c_out => CSA_carry_0_33_5);
FA_lbl_0_33_6: FA port map(in1 => b_and_a(653), in2 => b_and_a(684), c_in => b_and_a(715), sum => CSA_sum_0_33_6, c_out => CSA_carry_0_33_6);
FA_lbl_0_33_7: FA port map(in1 => b_and_a(746), in2 => b_and_a(777), c_in => b_and_a(808), sum => CSA_sum_0_33_7, c_out => CSA_carry_0_33_7);
FA_lbl_0_33_8: FA port map(in1 => b_and_a(839), in2 => b_and_a(870), c_in => b_and_a(901), sum => CSA_sum_0_33_8, c_out => CSA_carry_0_33_8);
FA_lbl_0_33_9: FA port map(in1 => b_and_a(932), in2 => b_and_a(963), c_in => b_and_a(994), sum => CSA_sum_0_33_9, c_out => CSA_carry_0_33_9);
FA_lbl_0_34_0: FA port map(in1 => b_and_a(127), in2 => b_and_a(158), c_in => b_and_a(189), sum => CSA_sum_0_34_0, c_out => CSA_carry_0_34_0);
FA_lbl_0_34_1: FA port map(in1 => b_and_a(220), in2 => b_and_a(251), c_in => b_and_a(282), sum => CSA_sum_0_34_1, c_out => CSA_carry_0_34_1);
FA_lbl_0_34_2: FA port map(in1 => b_and_a(313), in2 => b_and_a(344), c_in => b_and_a(375), sum => CSA_sum_0_34_2, c_out => CSA_carry_0_34_2);
FA_lbl_0_34_3: FA port map(in1 => b_and_a(406), in2 => b_and_a(437), c_in => b_and_a(468), sum => CSA_sum_0_34_3, c_out => CSA_carry_0_34_3);
FA_lbl_0_34_4: FA port map(in1 => b_and_a(499), in2 => b_and_a(530), c_in => b_and_a(561), sum => CSA_sum_0_34_4, c_out => CSA_carry_0_34_4);
FA_lbl_0_34_5: FA port map(in1 => b_and_a(592), in2 => b_and_a(623), c_in => b_and_a(654), sum => CSA_sum_0_34_5, c_out => CSA_carry_0_34_5);
FA_lbl_0_34_6: FA port map(in1 => b_and_a(685), in2 => b_and_a(716), c_in => b_and_a(747), sum => CSA_sum_0_34_6, c_out => CSA_carry_0_34_6);
FA_lbl_0_34_7: FA port map(in1 => b_and_a(778), in2 => b_and_a(809), c_in => b_and_a(840), sum => CSA_sum_0_34_7, c_out => CSA_carry_0_34_7);
FA_lbl_0_34_8: FA port map(in1 => b_and_a(871), in2 => b_and_a(902), c_in => b_and_a(933), sum => CSA_sum_0_34_8, c_out => CSA_carry_0_34_8);
FA_lbl_0_35_0: FA port map(in1 => b_and_a(159), in2 => b_and_a(190), c_in => b_and_a(221), sum => CSA_sum_0_35_0, c_out => CSA_carry_0_35_0);
FA_lbl_0_35_1: FA port map(in1 => b_and_a(252), in2 => b_and_a(283), c_in => b_and_a(314), sum => CSA_sum_0_35_1, c_out => CSA_carry_0_35_1);
FA_lbl_0_35_2: FA port map(in1 => b_and_a(345), in2 => b_and_a(376), c_in => b_and_a(407), sum => CSA_sum_0_35_2, c_out => CSA_carry_0_35_2);
FA_lbl_0_35_3: FA port map(in1 => b_and_a(438), in2 => b_and_a(469), c_in => b_and_a(500), sum => CSA_sum_0_35_3, c_out => CSA_carry_0_35_3);
FA_lbl_0_35_4: FA port map(in1 => b_and_a(531), in2 => b_and_a(562), c_in => b_and_a(593), sum => CSA_sum_0_35_4, c_out => CSA_carry_0_35_4);
FA_lbl_0_35_5: FA port map(in1 => b_and_a(624), in2 => b_and_a(655), c_in => b_and_a(686), sum => CSA_sum_0_35_5, c_out => CSA_carry_0_35_5);
FA_lbl_0_35_6: FA port map(in1 => b_and_a(717), in2 => b_and_a(748), c_in => b_and_a(779), sum => CSA_sum_0_35_6, c_out => CSA_carry_0_35_6);
FA_lbl_0_35_7: FA port map(in1 => b_and_a(810), in2 => b_and_a(841), c_in => b_and_a(872), sum => CSA_sum_0_35_7, c_out => CSA_carry_0_35_7);
FA_lbl_0_35_8: FA port map(in1 => b_and_a(903), in2 => b_and_a(934), c_in => b_and_a(965), sum => CSA_sum_0_35_8, c_out => CSA_carry_0_35_8);
FA_lbl_0_36_0: FA port map(in1 => b_and_a(191), in2 => b_and_a(222), c_in => b_and_a(253), sum => CSA_sum_0_36_0, c_out => CSA_carry_0_36_0);
FA_lbl_0_36_1: FA port map(in1 => b_and_a(284), in2 => b_and_a(315), c_in => b_and_a(346), sum => CSA_sum_0_36_1, c_out => CSA_carry_0_36_1);
FA_lbl_0_36_2: FA port map(in1 => b_and_a(377), in2 => b_and_a(408), c_in => b_and_a(439), sum => CSA_sum_0_36_2, c_out => CSA_carry_0_36_2);
FA_lbl_0_36_3: FA port map(in1 => b_and_a(470), in2 => b_and_a(501), c_in => b_and_a(532), sum => CSA_sum_0_36_3, c_out => CSA_carry_0_36_3);
FA_lbl_0_36_4: FA port map(in1 => b_and_a(563), in2 => b_and_a(594), c_in => b_and_a(625), sum => CSA_sum_0_36_4, c_out => CSA_carry_0_36_4);
FA_lbl_0_36_5: FA port map(in1 => b_and_a(656), in2 => b_and_a(687), c_in => b_and_a(718), sum => CSA_sum_0_36_5, c_out => CSA_carry_0_36_5);
FA_lbl_0_36_6: FA port map(in1 => b_and_a(749), in2 => b_and_a(780), c_in => b_and_a(811), sum => CSA_sum_0_36_6, c_out => CSA_carry_0_36_6);
FA_lbl_0_36_7: FA port map(in1 => b_and_a(842), in2 => b_and_a(873), c_in => b_and_a(904), sum => CSA_sum_0_36_7, c_out => CSA_carry_0_36_7);
FA_lbl_0_36_8: FA port map(in1 => b_and_a(935), in2 => b_and_a(966), c_in => b_and_a(997), sum => CSA_sum_0_36_8, c_out => CSA_carry_0_36_8);
FA_lbl_0_37_0: FA port map(in1 => b_and_a(223), in2 => b_and_a(254), c_in => b_and_a(285), sum => CSA_sum_0_37_0, c_out => CSA_carry_0_37_0);
FA_lbl_0_37_1: FA port map(in1 => b_and_a(316), in2 => b_and_a(347), c_in => b_and_a(378), sum => CSA_sum_0_37_1, c_out => CSA_carry_0_37_1);
FA_lbl_0_37_2: FA port map(in1 => b_and_a(409), in2 => b_and_a(440), c_in => b_and_a(471), sum => CSA_sum_0_37_2, c_out => CSA_carry_0_37_2);
FA_lbl_0_37_3: FA port map(in1 => b_and_a(502), in2 => b_and_a(533), c_in => b_and_a(564), sum => CSA_sum_0_37_3, c_out => CSA_carry_0_37_3);
FA_lbl_0_37_4: FA port map(in1 => b_and_a(595), in2 => b_and_a(626), c_in => b_and_a(657), sum => CSA_sum_0_37_4, c_out => CSA_carry_0_37_4);
FA_lbl_0_37_5: FA port map(in1 => b_and_a(688), in2 => b_and_a(719), c_in => b_and_a(750), sum => CSA_sum_0_37_5, c_out => CSA_carry_0_37_5);
FA_lbl_0_37_6: FA port map(in1 => b_and_a(781), in2 => b_and_a(812), c_in => b_and_a(843), sum => CSA_sum_0_37_6, c_out => CSA_carry_0_37_6);
FA_lbl_0_37_7: FA port map(in1 => b_and_a(874), in2 => b_and_a(905), c_in => b_and_a(936), sum => CSA_sum_0_37_7, c_out => CSA_carry_0_37_7);
FA_lbl_0_38_0: FA port map(in1 => b_and_a(255), in2 => b_and_a(286), c_in => b_and_a(317), sum => CSA_sum_0_38_0, c_out => CSA_carry_0_38_0);
FA_lbl_0_38_1: FA port map(in1 => b_and_a(348), in2 => b_and_a(379), c_in => b_and_a(410), sum => CSA_sum_0_38_1, c_out => CSA_carry_0_38_1);
FA_lbl_0_38_2: FA port map(in1 => b_and_a(441), in2 => b_and_a(472), c_in => b_and_a(503), sum => CSA_sum_0_38_2, c_out => CSA_carry_0_38_2);
FA_lbl_0_38_3: FA port map(in1 => b_and_a(534), in2 => b_and_a(565), c_in => b_and_a(596), sum => CSA_sum_0_38_3, c_out => CSA_carry_0_38_3);
FA_lbl_0_38_4: FA port map(in1 => b_and_a(627), in2 => b_and_a(658), c_in => b_and_a(689), sum => CSA_sum_0_38_4, c_out => CSA_carry_0_38_4);
FA_lbl_0_38_5: FA port map(in1 => b_and_a(720), in2 => b_and_a(751), c_in => b_and_a(782), sum => CSA_sum_0_38_5, c_out => CSA_carry_0_38_5);
FA_lbl_0_38_6: FA port map(in1 => b_and_a(813), in2 => b_and_a(844), c_in => b_and_a(875), sum => CSA_sum_0_38_6, c_out => CSA_carry_0_38_6);
FA_lbl_0_38_7: FA port map(in1 => b_and_a(906), in2 => b_and_a(937), c_in => b_and_a(968), sum => CSA_sum_0_38_7, c_out => CSA_carry_0_38_7);
FA_lbl_0_39_0: FA port map(in1 => b_and_a(287), in2 => b_and_a(318), c_in => b_and_a(349), sum => CSA_sum_0_39_0, c_out => CSA_carry_0_39_0);
FA_lbl_0_39_1: FA port map(in1 => b_and_a(380), in2 => b_and_a(411), c_in => b_and_a(442), sum => CSA_sum_0_39_1, c_out => CSA_carry_0_39_1);
FA_lbl_0_39_2: FA port map(in1 => b_and_a(473), in2 => b_and_a(504), c_in => b_and_a(535), sum => CSA_sum_0_39_2, c_out => CSA_carry_0_39_2);
FA_lbl_0_39_3: FA port map(in1 => b_and_a(566), in2 => b_and_a(597), c_in => b_and_a(628), sum => CSA_sum_0_39_3, c_out => CSA_carry_0_39_3);
FA_lbl_0_39_4: FA port map(in1 => b_and_a(659), in2 => b_and_a(690), c_in => b_and_a(721), sum => CSA_sum_0_39_4, c_out => CSA_carry_0_39_4);
FA_lbl_0_39_5: FA port map(in1 => b_and_a(752), in2 => b_and_a(783), c_in => b_and_a(814), sum => CSA_sum_0_39_5, c_out => CSA_carry_0_39_5);
FA_lbl_0_39_6: FA port map(in1 => b_and_a(845), in2 => b_and_a(876), c_in => b_and_a(907), sum => CSA_sum_0_39_6, c_out => CSA_carry_0_39_6);
FA_lbl_0_39_7: FA port map(in1 => b_and_a(938), in2 => b_and_a(969), c_in => b_and_a(1000), sum => CSA_sum_0_39_7, c_out => CSA_carry_0_39_7);
FA_lbl_0_40_0: FA port map(in1 => b_and_a(319), in2 => b_and_a(350), c_in => b_and_a(381), sum => CSA_sum_0_40_0, c_out => CSA_carry_0_40_0);
FA_lbl_0_40_1: FA port map(in1 => b_and_a(412), in2 => b_and_a(443), c_in => b_and_a(474), sum => CSA_sum_0_40_1, c_out => CSA_carry_0_40_1);
FA_lbl_0_40_2: FA port map(in1 => b_and_a(505), in2 => b_and_a(536), c_in => b_and_a(567), sum => CSA_sum_0_40_2, c_out => CSA_carry_0_40_2);
FA_lbl_0_40_3: FA port map(in1 => b_and_a(598), in2 => b_and_a(629), c_in => b_and_a(660), sum => CSA_sum_0_40_3, c_out => CSA_carry_0_40_3);
FA_lbl_0_40_4: FA port map(in1 => b_and_a(691), in2 => b_and_a(722), c_in => b_and_a(753), sum => CSA_sum_0_40_4, c_out => CSA_carry_0_40_4);
FA_lbl_0_40_5: FA port map(in1 => b_and_a(784), in2 => b_and_a(815), c_in => b_and_a(846), sum => CSA_sum_0_40_5, c_out => CSA_carry_0_40_5);
FA_lbl_0_40_6: FA port map(in1 => b_and_a(877), in2 => b_and_a(908), c_in => b_and_a(939), sum => CSA_sum_0_40_6, c_out => CSA_carry_0_40_6);
FA_lbl_0_41_0: FA port map(in1 => b_and_a(351), in2 => b_and_a(382), c_in => b_and_a(413), sum => CSA_sum_0_41_0, c_out => CSA_carry_0_41_0);
FA_lbl_0_41_1: FA port map(in1 => b_and_a(444), in2 => b_and_a(475), c_in => b_and_a(506), sum => CSA_sum_0_41_1, c_out => CSA_carry_0_41_1);
FA_lbl_0_41_2: FA port map(in1 => b_and_a(537), in2 => b_and_a(568), c_in => b_and_a(599), sum => CSA_sum_0_41_2, c_out => CSA_carry_0_41_2);
FA_lbl_0_41_3: FA port map(in1 => b_and_a(630), in2 => b_and_a(661), c_in => b_and_a(692), sum => CSA_sum_0_41_3, c_out => CSA_carry_0_41_3);
FA_lbl_0_41_4: FA port map(in1 => b_and_a(723), in2 => b_and_a(754), c_in => b_and_a(785), sum => CSA_sum_0_41_4, c_out => CSA_carry_0_41_4);
FA_lbl_0_41_5: FA port map(in1 => b_and_a(816), in2 => b_and_a(847), c_in => b_and_a(878), sum => CSA_sum_0_41_5, c_out => CSA_carry_0_41_5);
FA_lbl_0_41_6: FA port map(in1 => b_and_a(909), in2 => b_and_a(940), c_in => b_and_a(971), sum => CSA_sum_0_41_6, c_out => CSA_carry_0_41_6);
FA_lbl_0_42_0: FA port map(in1 => b_and_a(383), in2 => b_and_a(414), c_in => b_and_a(445), sum => CSA_sum_0_42_0, c_out => CSA_carry_0_42_0);
FA_lbl_0_42_1: FA port map(in1 => b_and_a(476), in2 => b_and_a(507), c_in => b_and_a(538), sum => CSA_sum_0_42_1, c_out => CSA_carry_0_42_1);
FA_lbl_0_42_2: FA port map(in1 => b_and_a(569), in2 => b_and_a(600), c_in => b_and_a(631), sum => CSA_sum_0_42_2, c_out => CSA_carry_0_42_2);
FA_lbl_0_42_3: FA port map(in1 => b_and_a(662), in2 => b_and_a(693), c_in => b_and_a(724), sum => CSA_sum_0_42_3, c_out => CSA_carry_0_42_3);
FA_lbl_0_42_4: FA port map(in1 => b_and_a(755), in2 => b_and_a(786), c_in => b_and_a(817), sum => CSA_sum_0_42_4, c_out => CSA_carry_0_42_4);
FA_lbl_0_42_5: FA port map(in1 => b_and_a(848), in2 => b_and_a(879), c_in => b_and_a(910), sum => CSA_sum_0_42_5, c_out => CSA_carry_0_42_5);
FA_lbl_0_42_6: FA port map(in1 => b_and_a(941), in2 => b_and_a(972), c_in => b_and_a(1003), sum => CSA_sum_0_42_6, c_out => CSA_carry_0_42_6);
FA_lbl_0_43_0: FA port map(in1 => b_and_a(415), in2 => b_and_a(446), c_in => b_and_a(477), sum => CSA_sum_0_43_0, c_out => CSA_carry_0_43_0);
FA_lbl_0_43_1: FA port map(in1 => b_and_a(508), in2 => b_and_a(539), c_in => b_and_a(570), sum => CSA_sum_0_43_1, c_out => CSA_carry_0_43_1);
FA_lbl_0_43_2: FA port map(in1 => b_and_a(601), in2 => b_and_a(632), c_in => b_and_a(663), sum => CSA_sum_0_43_2, c_out => CSA_carry_0_43_2);
FA_lbl_0_43_3: FA port map(in1 => b_and_a(694), in2 => b_and_a(725), c_in => b_and_a(756), sum => CSA_sum_0_43_3, c_out => CSA_carry_0_43_3);
FA_lbl_0_43_4: FA port map(in1 => b_and_a(787), in2 => b_and_a(818), c_in => b_and_a(849), sum => CSA_sum_0_43_4, c_out => CSA_carry_0_43_4);
FA_lbl_0_43_5: FA port map(in1 => b_and_a(880), in2 => b_and_a(911), c_in => b_and_a(942), sum => CSA_sum_0_43_5, c_out => CSA_carry_0_43_5);
FA_lbl_0_44_0: FA port map(in1 => b_and_a(447), in2 => b_and_a(478), c_in => b_and_a(509), sum => CSA_sum_0_44_0, c_out => CSA_carry_0_44_0);
FA_lbl_0_44_1: FA port map(in1 => b_and_a(540), in2 => b_and_a(571), c_in => b_and_a(602), sum => CSA_sum_0_44_1, c_out => CSA_carry_0_44_1);
FA_lbl_0_44_2: FA port map(in1 => b_and_a(633), in2 => b_and_a(664), c_in => b_and_a(695), sum => CSA_sum_0_44_2, c_out => CSA_carry_0_44_2);
FA_lbl_0_44_3: FA port map(in1 => b_and_a(726), in2 => b_and_a(757), c_in => b_and_a(788), sum => CSA_sum_0_44_3, c_out => CSA_carry_0_44_3);
FA_lbl_0_44_4: FA port map(in1 => b_and_a(819), in2 => b_and_a(850), c_in => b_and_a(881), sum => CSA_sum_0_44_4, c_out => CSA_carry_0_44_4);
FA_lbl_0_44_5: FA port map(in1 => b_and_a(912), in2 => b_and_a(943), c_in => b_and_a(974), sum => CSA_sum_0_44_5, c_out => CSA_carry_0_44_5);
FA_lbl_0_45_0: FA port map(in1 => b_and_a(479), in2 => b_and_a(510), c_in => b_and_a(541), sum => CSA_sum_0_45_0, c_out => CSA_carry_0_45_0);
FA_lbl_0_45_1: FA port map(in1 => b_and_a(572), in2 => b_and_a(603), c_in => b_and_a(634), sum => CSA_sum_0_45_1, c_out => CSA_carry_0_45_1);
FA_lbl_0_45_2: FA port map(in1 => b_and_a(665), in2 => b_and_a(696), c_in => b_and_a(727), sum => CSA_sum_0_45_2, c_out => CSA_carry_0_45_2);
FA_lbl_0_45_3: FA port map(in1 => b_and_a(758), in2 => b_and_a(789), c_in => b_and_a(820), sum => CSA_sum_0_45_3, c_out => CSA_carry_0_45_3);
FA_lbl_0_45_4: FA port map(in1 => b_and_a(851), in2 => b_and_a(882), c_in => b_and_a(913), sum => CSA_sum_0_45_4, c_out => CSA_carry_0_45_4);
FA_lbl_0_45_5: FA port map(in1 => b_and_a(944), in2 => b_and_a(975), c_in => b_and_a(1006), sum => CSA_sum_0_45_5, c_out => CSA_carry_0_45_5);
FA_lbl_0_46_0: FA port map(in1 => b_and_a(511), in2 => b_and_a(542), c_in => b_and_a(573), sum => CSA_sum_0_46_0, c_out => CSA_carry_0_46_0);
FA_lbl_0_46_1: FA port map(in1 => b_and_a(604), in2 => b_and_a(635), c_in => b_and_a(666), sum => CSA_sum_0_46_1, c_out => CSA_carry_0_46_1);
FA_lbl_0_46_2: FA port map(in1 => b_and_a(697), in2 => b_and_a(728), c_in => b_and_a(759), sum => CSA_sum_0_46_2, c_out => CSA_carry_0_46_2);
FA_lbl_0_46_3: FA port map(in1 => b_and_a(790), in2 => b_and_a(821), c_in => b_and_a(852), sum => CSA_sum_0_46_3, c_out => CSA_carry_0_46_3);
FA_lbl_0_46_4: FA port map(in1 => b_and_a(883), in2 => b_and_a(914), c_in => b_and_a(945), sum => CSA_sum_0_46_4, c_out => CSA_carry_0_46_4);
FA_lbl_0_47_0: FA port map(in1 => b_and_a(543), in2 => b_and_a(574), c_in => b_and_a(605), sum => CSA_sum_0_47_0, c_out => CSA_carry_0_47_0);
FA_lbl_0_47_1: FA port map(in1 => b_and_a(636), in2 => b_and_a(667), c_in => b_and_a(698), sum => CSA_sum_0_47_1, c_out => CSA_carry_0_47_1);
FA_lbl_0_47_2: FA port map(in1 => b_and_a(729), in2 => b_and_a(760), c_in => b_and_a(791), sum => CSA_sum_0_47_2, c_out => CSA_carry_0_47_2);
FA_lbl_0_47_3: FA port map(in1 => b_and_a(822), in2 => b_and_a(853), c_in => b_and_a(884), sum => CSA_sum_0_47_3, c_out => CSA_carry_0_47_3);
FA_lbl_0_47_4: FA port map(in1 => b_and_a(915), in2 => b_and_a(946), c_in => b_and_a(977), sum => CSA_sum_0_47_4, c_out => CSA_carry_0_47_4);
FA_lbl_0_48_0: FA port map(in1 => b_and_a(575), in2 => b_and_a(606), c_in => b_and_a(637), sum => CSA_sum_0_48_0, c_out => CSA_carry_0_48_0);
FA_lbl_0_48_1: FA port map(in1 => b_and_a(668), in2 => b_and_a(699), c_in => b_and_a(730), sum => CSA_sum_0_48_1, c_out => CSA_carry_0_48_1);
FA_lbl_0_48_2: FA port map(in1 => b_and_a(761), in2 => b_and_a(792), c_in => b_and_a(823), sum => CSA_sum_0_48_2, c_out => CSA_carry_0_48_2);
FA_lbl_0_48_3: FA port map(in1 => b_and_a(854), in2 => b_and_a(885), c_in => b_and_a(916), sum => CSA_sum_0_48_3, c_out => CSA_carry_0_48_3);
FA_lbl_0_48_4: FA port map(in1 => b_and_a(947), in2 => b_and_a(978), c_in => b_and_a(1009), sum => CSA_sum_0_48_4, c_out => CSA_carry_0_48_4);
FA_lbl_0_49_0: FA port map(in1 => b_and_a(607), in2 => b_and_a(638), c_in => b_and_a(669), sum => CSA_sum_0_49_0, c_out => CSA_carry_0_49_0);
FA_lbl_0_49_1: FA port map(in1 => b_and_a(700), in2 => b_and_a(731), c_in => b_and_a(762), sum => CSA_sum_0_49_1, c_out => CSA_carry_0_49_1);
FA_lbl_0_49_2: FA port map(in1 => b_and_a(793), in2 => b_and_a(824), c_in => b_and_a(855), sum => CSA_sum_0_49_2, c_out => CSA_carry_0_49_2);
FA_lbl_0_49_3: FA port map(in1 => b_and_a(886), in2 => b_and_a(917), c_in => b_and_a(948), sum => CSA_sum_0_49_3, c_out => CSA_carry_0_49_3);
FA_lbl_0_50_0: FA port map(in1 => b_and_a(639), in2 => b_and_a(670), c_in => b_and_a(701), sum => CSA_sum_0_50_0, c_out => CSA_carry_0_50_0);
FA_lbl_0_50_1: FA port map(in1 => b_and_a(732), in2 => b_and_a(763), c_in => b_and_a(794), sum => CSA_sum_0_50_1, c_out => CSA_carry_0_50_1);
FA_lbl_0_50_2: FA port map(in1 => b_and_a(825), in2 => b_and_a(856), c_in => b_and_a(887), sum => CSA_sum_0_50_2, c_out => CSA_carry_0_50_2);
FA_lbl_0_50_3: FA port map(in1 => b_and_a(918), in2 => b_and_a(949), c_in => b_and_a(980), sum => CSA_sum_0_50_3, c_out => CSA_carry_0_50_3);
FA_lbl_0_51_0: FA port map(in1 => b_and_a(671), in2 => b_and_a(702), c_in => b_and_a(733), sum => CSA_sum_0_51_0, c_out => CSA_carry_0_51_0);
FA_lbl_0_51_1: FA port map(in1 => b_and_a(764), in2 => b_and_a(795), c_in => b_and_a(826), sum => CSA_sum_0_51_1, c_out => CSA_carry_0_51_1);
FA_lbl_0_51_2: FA port map(in1 => b_and_a(857), in2 => b_and_a(888), c_in => b_and_a(919), sum => CSA_sum_0_51_2, c_out => CSA_carry_0_51_2);
FA_lbl_0_51_3: FA port map(in1 => b_and_a(950), in2 => b_and_a(981), c_in => b_and_a(1012), sum => CSA_sum_0_51_3, c_out => CSA_carry_0_51_3);
FA_lbl_0_52_0: FA port map(in1 => b_and_a(703), in2 => b_and_a(734), c_in => b_and_a(765), sum => CSA_sum_0_52_0, c_out => CSA_carry_0_52_0);
FA_lbl_0_52_1: FA port map(in1 => b_and_a(796), in2 => b_and_a(827), c_in => b_and_a(858), sum => CSA_sum_0_52_1, c_out => CSA_carry_0_52_1);
FA_lbl_0_52_2: FA port map(in1 => b_and_a(889), in2 => b_and_a(920), c_in => b_and_a(951), sum => CSA_sum_0_52_2, c_out => CSA_carry_0_52_2);
FA_lbl_0_53_0: FA port map(in1 => b_and_a(735), in2 => b_and_a(766), c_in => b_and_a(797), sum => CSA_sum_0_53_0, c_out => CSA_carry_0_53_0);
FA_lbl_0_53_1: FA port map(in1 => b_and_a(828), in2 => b_and_a(859), c_in => b_and_a(890), sum => CSA_sum_0_53_1, c_out => CSA_carry_0_53_1);
FA_lbl_0_53_2: FA port map(in1 => b_and_a(921), in2 => b_and_a(952), c_in => b_and_a(983), sum => CSA_sum_0_53_2, c_out => CSA_carry_0_53_2);
FA_lbl_0_54_0: FA port map(in1 => b_and_a(767), in2 => b_and_a(798), c_in => b_and_a(829), sum => CSA_sum_0_54_0, c_out => CSA_carry_0_54_0);
FA_lbl_0_54_1: FA port map(in1 => b_and_a(860), in2 => b_and_a(891), c_in => b_and_a(922), sum => CSA_sum_0_54_1, c_out => CSA_carry_0_54_1);
FA_lbl_0_54_2: FA port map(in1 => b_and_a(953), in2 => b_and_a(984), c_in => b_and_a(1015), sum => CSA_sum_0_54_2, c_out => CSA_carry_0_54_2);
FA_lbl_0_55_0: FA port map(in1 => b_and_a(799), in2 => b_and_a(830), c_in => b_and_a(861), sum => CSA_sum_0_55_0, c_out => CSA_carry_0_55_0);
FA_lbl_0_55_1: FA port map(in1 => b_and_a(892), in2 => b_and_a(923), c_in => b_and_a(954), sum => CSA_sum_0_55_1, c_out => CSA_carry_0_55_1);
FA_lbl_0_56_0: FA port map(in1 => b_and_a(831), in2 => b_and_a(862), c_in => b_and_a(893), sum => CSA_sum_0_56_0, c_out => CSA_carry_0_56_0);
FA_lbl_0_56_1: FA port map(in1 => b_and_a(924), in2 => b_and_a(955), c_in => b_and_a(986), sum => CSA_sum_0_56_1, c_out => CSA_carry_0_56_1);
FA_lbl_0_57_0: FA port map(in1 => b_and_a(863), in2 => b_and_a(894), c_in => b_and_a(925), sum => CSA_sum_0_57_0, c_out => CSA_carry_0_57_0);
FA_lbl_0_57_1: FA port map(in1 => b_and_a(956), in2 => b_and_a(987), c_in => b_and_a(1018), sum => CSA_sum_0_57_1, c_out => CSA_carry_0_57_1);
FA_lbl_0_58_0: FA port map(in1 => b_and_a(895), in2 => b_and_a(926), c_in => b_and_a(957), sum => CSA_sum_0_58_0, c_out => CSA_carry_0_58_0);
FA_lbl_0_59_0: FA port map(in1 => b_and_a(927), in2 => b_and_a(958), c_in => b_and_a(989), sum => CSA_sum_0_59_0, c_out => CSA_carry_0_59_0);
FA_lbl_0_60_0: FA port map(in1 => b_and_a(959), in2 => b_and_a(990), c_in => b_and_a(1021), sum => CSA_sum_0_60_0, c_out => CSA_carry_0_60_0);
FA_lbl_1_3_0: FA port map(in1 => b_and_a(96), in2 => CSA_sum_0_3_0, c_in => CSA_carry_0_2_0, sum => CSA_sum_1_3_0, c_out => CSA_carry_1_3_0);
FA_lbl_1_4_0: FA port map(in1 => b_and_a(97), in2 => b_and_a(128), c_in => CSA_sum_0_4_0, sum => CSA_sum_1_4_0, c_out => CSA_carry_1_4_0);
FA_lbl_1_5_0: FA port map(in1 => CSA_sum_0_5_1, in2 => CSA_sum_0_5_0, c_in => CSA_carry_0_4_0, sum => CSA_sum_1_5_0, c_out => CSA_carry_1_5_0);
FA_lbl_1_6_0: FA port map(in1 => b_and_a(192), in2 => CSA_sum_0_6_1, c_in => CSA_sum_0_6_0, sum => CSA_sum_1_6_0, c_out => CSA_carry_1_6_0);
FA_lbl_1_7_0: FA port map(in1 => b_and_a(193), in2 => b_and_a(224), c_in => CSA_sum_0_7_1, sum => CSA_sum_1_7_0, c_out => CSA_carry_1_7_0);
FA_lbl_1_7_1: FA port map(in1 => CSA_sum_0_7_0, in2 => CSA_carry_0_6_1, c_in => CSA_carry_0_6_0, sum => CSA_sum_1_7_1, c_out => CSA_carry_1_7_1);
FA_lbl_1_8_0: FA port map(in1 => CSA_sum_0_8_2, in2 => CSA_sum_0_8_1, c_in => CSA_sum_0_8_0, sum => CSA_sum_1_8_0, c_out => CSA_carry_1_8_0);
FA_lbl_1_9_0: FA port map(in1 => b_and_a(288), in2 => CSA_sum_0_9_2, c_in => CSA_sum_0_9_1, sum => CSA_sum_1_9_0, c_out => CSA_carry_1_9_0);
FA_lbl_1_9_1: FA port map(in1 => CSA_sum_0_9_0, in2 => CSA_carry_0_8_2, c_in => CSA_carry_0_8_1, sum => CSA_sum_1_9_1, c_out => CSA_carry_1_9_1);
FA_lbl_1_10_0: FA port map(in1 => b_and_a(289), in2 => b_and_a(320), c_in => CSA_sum_0_10_2, sum => CSA_sum_1_10_0, c_out => CSA_carry_1_10_0);
FA_lbl_1_10_1: FA port map(in1 => CSA_sum_0_10_1, in2 => CSA_sum_0_10_0, c_in => CSA_carry_0_9_2, sum => CSA_sum_1_10_1, c_out => CSA_carry_1_10_1);
FA_lbl_1_11_0: FA port map(in1 => CSA_sum_0_11_3, in2 => CSA_sum_0_11_2, c_in => CSA_sum_0_11_1, sum => CSA_sum_1_11_0, c_out => CSA_carry_1_11_0);
FA_lbl_1_11_1: FA port map(in1 => CSA_sum_0_11_0, in2 => CSA_carry_0_10_2, c_in => CSA_carry_0_10_1, sum => CSA_sum_1_11_1, c_out => CSA_carry_1_11_1);
FA_lbl_1_12_0: FA port map(in1 => b_and_a(384), in2 => CSA_sum_0_12_3, c_in => CSA_sum_0_12_2, sum => CSA_sum_1_12_0, c_out => CSA_carry_1_12_0);
FA_lbl_1_12_1: FA port map(in1 => CSA_sum_0_12_1, in2 => CSA_sum_0_12_0, c_in => CSA_carry_0_11_3, sum => CSA_sum_1_12_1, c_out => CSA_carry_1_12_1);
FA_lbl_1_12_2: FA port map(in1 => CSA_carry_0_11_2, in2 => CSA_carry_0_11_1, c_in => CSA_carry_0_11_0, sum => CSA_sum_1_12_2, c_out => CSA_carry_1_12_2);
FA_lbl_1_13_0: FA port map(in1 => b_and_a(385), in2 => b_and_a(416), c_in => CSA_sum_0_13_3, sum => CSA_sum_1_13_0, c_out => CSA_carry_1_13_0);
FA_lbl_1_13_1: FA port map(in1 => CSA_sum_0_13_2, in2 => CSA_sum_0_13_1, c_in => CSA_sum_0_13_0, sum => CSA_sum_1_13_1, c_out => CSA_carry_1_13_1);
FA_lbl_1_13_2: FA port map(in1 => CSA_carry_0_12_3, in2 => CSA_carry_0_12_2, c_in => CSA_carry_0_12_1, sum => CSA_sum_1_13_2, c_out => CSA_carry_1_13_2);
FA_lbl_1_14_0: FA port map(in1 => CSA_sum_0_14_4, in2 => CSA_sum_0_14_3, c_in => CSA_sum_0_14_2, sum => CSA_sum_1_14_0, c_out => CSA_carry_1_14_0);
FA_lbl_1_14_1: FA port map(in1 => CSA_sum_0_14_1, in2 => CSA_sum_0_14_0, c_in => CSA_carry_0_13_3, sum => CSA_sum_1_14_1, c_out => CSA_carry_1_14_1);
FA_lbl_1_14_2: FA port map(in1 => CSA_carry_0_13_2, in2 => CSA_carry_0_13_1, c_in => CSA_carry_0_13_0, sum => CSA_sum_1_14_2, c_out => CSA_carry_1_14_2);
FA_lbl_1_15_0: FA port map(in1 => b_and_a(480), in2 => CSA_sum_0_15_4, c_in => CSA_sum_0_15_3, sum => CSA_sum_1_15_0, c_out => CSA_carry_1_15_0);
FA_lbl_1_15_1: FA port map(in1 => CSA_sum_0_15_2, in2 => CSA_sum_0_15_1, c_in => CSA_sum_0_15_0, sum => CSA_sum_1_15_1, c_out => CSA_carry_1_15_1);
FA_lbl_1_15_2: FA port map(in1 => CSA_carry_0_14_4, in2 => CSA_carry_0_14_3, c_in => CSA_carry_0_14_2, sum => CSA_sum_1_15_2, c_out => CSA_carry_1_15_2);
FA_lbl_1_16_0: FA port map(in1 => b_and_a(481), in2 => b_and_a(512), c_in => CSA_sum_0_16_4, sum => CSA_sum_1_16_0, c_out => CSA_carry_1_16_0);
FA_lbl_1_16_1: FA port map(in1 => CSA_sum_0_16_3, in2 => CSA_sum_0_16_2, c_in => CSA_sum_0_16_1, sum => CSA_sum_1_16_1, c_out => CSA_carry_1_16_1);
FA_lbl_1_16_2: FA port map(in1 => CSA_sum_0_16_0, in2 => CSA_carry_0_15_4, c_in => CSA_carry_0_15_3, sum => CSA_sum_1_16_2, c_out => CSA_carry_1_16_2);
FA_lbl_1_16_3: FA port map(in1 => CSA_carry_0_15_2, in2 => CSA_carry_0_15_1, c_in => CSA_carry_0_15_0, sum => CSA_sum_1_16_3, c_out => CSA_carry_1_16_3);
FA_lbl_1_17_0: FA port map(in1 => CSA_sum_0_17_5, in2 => CSA_sum_0_17_4, c_in => CSA_sum_0_17_3, sum => CSA_sum_1_17_0, c_out => CSA_carry_1_17_0);
FA_lbl_1_17_1: FA port map(in1 => CSA_sum_0_17_2, in2 => CSA_sum_0_17_1, c_in => CSA_sum_0_17_0, sum => CSA_sum_1_17_1, c_out => CSA_carry_1_17_1);
FA_lbl_1_17_2: FA port map(in1 => CSA_carry_0_16_4, in2 => CSA_carry_0_16_3, c_in => CSA_carry_0_16_2, sum => CSA_sum_1_17_2, c_out => CSA_carry_1_17_2);
FA_lbl_1_18_0: FA port map(in1 => b_and_a(576), in2 => CSA_sum_0_18_5, c_in => CSA_sum_0_18_4, sum => CSA_sum_1_18_0, c_out => CSA_carry_1_18_0);
FA_lbl_1_18_1: FA port map(in1 => CSA_sum_0_18_3, in2 => CSA_sum_0_18_2, c_in => CSA_sum_0_18_1, sum => CSA_sum_1_18_1, c_out => CSA_carry_1_18_1);
FA_lbl_1_18_2: FA port map(in1 => CSA_sum_0_18_0, in2 => CSA_carry_0_17_5, c_in => CSA_carry_0_17_4, sum => CSA_sum_1_18_2, c_out => CSA_carry_1_18_2);
FA_lbl_1_18_3: FA port map(in1 => CSA_carry_0_17_3, in2 => CSA_carry_0_17_2, c_in => CSA_carry_0_17_1, sum => CSA_sum_1_18_3, c_out => CSA_carry_1_18_3);
FA_lbl_1_19_0: FA port map(in1 => b_and_a(577), in2 => b_and_a(608), c_in => CSA_sum_0_19_5, sum => CSA_sum_1_19_0, c_out => CSA_carry_1_19_0);
FA_lbl_1_19_1: FA port map(in1 => CSA_sum_0_19_4, in2 => CSA_sum_0_19_3, c_in => CSA_sum_0_19_2, sum => CSA_sum_1_19_1, c_out => CSA_carry_1_19_1);
FA_lbl_1_19_2: FA port map(in1 => CSA_sum_0_19_1, in2 => CSA_sum_0_19_0, c_in => CSA_carry_0_18_5, sum => CSA_sum_1_19_2, c_out => CSA_carry_1_19_2);
FA_lbl_1_19_3: FA port map(in1 => CSA_carry_0_18_4, in2 => CSA_carry_0_18_3, c_in => CSA_carry_0_18_2, sum => CSA_sum_1_19_3, c_out => CSA_carry_1_19_3);
FA_lbl_1_20_0: FA port map(in1 => CSA_sum_0_20_6, in2 => CSA_sum_0_20_5, c_in => CSA_sum_0_20_4, sum => CSA_sum_1_20_0, c_out => CSA_carry_1_20_0);
FA_lbl_1_20_1: FA port map(in1 => CSA_sum_0_20_3, in2 => CSA_sum_0_20_2, c_in => CSA_sum_0_20_1, sum => CSA_sum_1_20_1, c_out => CSA_carry_1_20_1);
FA_lbl_1_20_2: FA port map(in1 => CSA_sum_0_20_0, in2 => CSA_carry_0_19_5, c_in => CSA_carry_0_19_4, sum => CSA_sum_1_20_2, c_out => CSA_carry_1_20_2);
FA_lbl_1_20_3: FA port map(in1 => CSA_carry_0_19_3, in2 => CSA_carry_0_19_2, c_in => CSA_carry_0_19_1, sum => CSA_sum_1_20_3, c_out => CSA_carry_1_20_3);
FA_lbl_1_21_0: FA port map(in1 => b_and_a(672), in2 => CSA_sum_0_21_6, c_in => CSA_sum_0_21_5, sum => CSA_sum_1_21_0, c_out => CSA_carry_1_21_0);
FA_lbl_1_21_1: FA port map(in1 => CSA_sum_0_21_4, in2 => CSA_sum_0_21_3, c_in => CSA_sum_0_21_2, sum => CSA_sum_1_21_1, c_out => CSA_carry_1_21_1);
FA_lbl_1_21_2: FA port map(in1 => CSA_sum_0_21_1, in2 => CSA_sum_0_21_0, c_in => CSA_carry_0_20_6, sum => CSA_sum_1_21_2, c_out => CSA_carry_1_21_2);
FA_lbl_1_21_3: FA port map(in1 => CSA_carry_0_20_5, in2 => CSA_carry_0_20_4, c_in => CSA_carry_0_20_3, sum => CSA_sum_1_21_3, c_out => CSA_carry_1_21_3);
FA_lbl_1_21_4: FA port map(in1 => CSA_carry_0_20_2, in2 => CSA_carry_0_20_1, c_in => CSA_carry_0_20_0, sum => CSA_sum_1_21_4, c_out => CSA_carry_1_21_4);
FA_lbl_1_22_0: FA port map(in1 => b_and_a(673), in2 => b_and_a(704), c_in => CSA_sum_0_22_6, sum => CSA_sum_1_22_0, c_out => CSA_carry_1_22_0);
FA_lbl_1_22_1: FA port map(in1 => CSA_sum_0_22_5, in2 => CSA_sum_0_22_4, c_in => CSA_sum_0_22_3, sum => CSA_sum_1_22_1, c_out => CSA_carry_1_22_1);
FA_lbl_1_22_2: FA port map(in1 => CSA_sum_0_22_2, in2 => CSA_sum_0_22_1, c_in => CSA_sum_0_22_0, sum => CSA_sum_1_22_2, c_out => CSA_carry_1_22_2);
FA_lbl_1_22_3: FA port map(in1 => CSA_carry_0_21_6, in2 => CSA_carry_0_21_5, c_in => CSA_carry_0_21_4, sum => CSA_sum_1_22_3, c_out => CSA_carry_1_22_3);
FA_lbl_1_22_4: FA port map(in1 => CSA_carry_0_21_3, in2 => CSA_carry_0_21_2, c_in => CSA_carry_0_21_1, sum => CSA_sum_1_22_4, c_out => CSA_carry_1_22_4);
FA_lbl_1_23_0: FA port map(in1 => CSA_sum_0_23_7, in2 => CSA_sum_0_23_6, c_in => CSA_sum_0_23_5, sum => CSA_sum_1_23_0, c_out => CSA_carry_1_23_0);
FA_lbl_1_23_1: FA port map(in1 => CSA_sum_0_23_4, in2 => CSA_sum_0_23_3, c_in => CSA_sum_0_23_2, sum => CSA_sum_1_23_1, c_out => CSA_carry_1_23_1);
FA_lbl_1_23_2: FA port map(in1 => CSA_sum_0_23_1, in2 => CSA_sum_0_23_0, c_in => CSA_carry_0_22_6, sum => CSA_sum_1_23_2, c_out => CSA_carry_1_23_2);
FA_lbl_1_23_3: FA port map(in1 => CSA_carry_0_22_5, in2 => CSA_carry_0_22_4, c_in => CSA_carry_0_22_3, sum => CSA_sum_1_23_3, c_out => CSA_carry_1_23_3);
FA_lbl_1_23_4: FA port map(in1 => CSA_carry_0_22_2, in2 => CSA_carry_0_22_1, c_in => CSA_carry_0_22_0, sum => CSA_sum_1_23_4, c_out => CSA_carry_1_23_4);
FA_lbl_1_24_0: FA port map(in1 => b_and_a(768), in2 => CSA_sum_0_24_7, c_in => CSA_sum_0_24_6, sum => CSA_sum_1_24_0, c_out => CSA_carry_1_24_0);
FA_lbl_1_24_1: FA port map(in1 => CSA_sum_0_24_5, in2 => CSA_sum_0_24_4, c_in => CSA_sum_0_24_3, sum => CSA_sum_1_24_1, c_out => CSA_carry_1_24_1);
FA_lbl_1_24_2: FA port map(in1 => CSA_sum_0_24_2, in2 => CSA_sum_0_24_1, c_in => CSA_sum_0_24_0, sum => CSA_sum_1_24_2, c_out => CSA_carry_1_24_2);
FA_lbl_1_24_3: FA port map(in1 => CSA_carry_0_23_7, in2 => CSA_carry_0_23_6, c_in => CSA_carry_0_23_5, sum => CSA_sum_1_24_3, c_out => CSA_carry_1_24_3);
FA_lbl_1_24_4: FA port map(in1 => CSA_carry_0_23_4, in2 => CSA_carry_0_23_3, c_in => CSA_carry_0_23_2, sum => CSA_sum_1_24_4, c_out => CSA_carry_1_24_4);
FA_lbl_1_25_0: FA port map(in1 => b_and_a(769), in2 => b_and_a(800), c_in => CSA_sum_0_25_7, sum => CSA_sum_1_25_0, c_out => CSA_carry_1_25_0);
FA_lbl_1_25_1: FA port map(in1 => CSA_sum_0_25_6, in2 => CSA_sum_0_25_5, c_in => CSA_sum_0_25_4, sum => CSA_sum_1_25_1, c_out => CSA_carry_1_25_1);
FA_lbl_1_25_2: FA port map(in1 => CSA_sum_0_25_3, in2 => CSA_sum_0_25_2, c_in => CSA_sum_0_25_1, sum => CSA_sum_1_25_2, c_out => CSA_carry_1_25_2);
FA_lbl_1_25_3: FA port map(in1 => CSA_sum_0_25_0, in2 => CSA_carry_0_24_7, c_in => CSA_carry_0_24_6, sum => CSA_sum_1_25_3, c_out => CSA_carry_1_25_3);
FA_lbl_1_25_4: FA port map(in1 => CSA_carry_0_24_5, in2 => CSA_carry_0_24_4, c_in => CSA_carry_0_24_3, sum => CSA_sum_1_25_4, c_out => CSA_carry_1_25_4);
FA_lbl_1_25_5: FA port map(in1 => CSA_carry_0_24_2, in2 => CSA_carry_0_24_1, c_in => CSA_carry_0_24_0, sum => CSA_sum_1_25_5, c_out => CSA_carry_1_25_5);
FA_lbl_1_26_0: FA port map(in1 => CSA_sum_0_26_8, in2 => CSA_sum_0_26_7, c_in => CSA_sum_0_26_6, sum => CSA_sum_1_26_0, c_out => CSA_carry_1_26_0);
FA_lbl_1_26_1: FA port map(in1 => CSA_sum_0_26_5, in2 => CSA_sum_0_26_4, c_in => CSA_sum_0_26_3, sum => CSA_sum_1_26_1, c_out => CSA_carry_1_26_1);
FA_lbl_1_26_2: FA port map(in1 => CSA_sum_0_26_2, in2 => CSA_sum_0_26_1, c_in => CSA_sum_0_26_0, sum => CSA_sum_1_26_2, c_out => CSA_carry_1_26_2);
FA_lbl_1_26_3: FA port map(in1 => CSA_carry_0_25_7, in2 => CSA_carry_0_25_6, c_in => CSA_carry_0_25_5, sum => CSA_sum_1_26_3, c_out => CSA_carry_1_26_3);
FA_lbl_1_26_4: FA port map(in1 => CSA_carry_0_25_4, in2 => CSA_carry_0_25_3, c_in => CSA_carry_0_25_2, sum => CSA_sum_1_26_4, c_out => CSA_carry_1_26_4);
FA_lbl_1_27_0: FA port map(in1 => b_and_a(864), in2 => CSA_sum_0_27_8, c_in => CSA_sum_0_27_7, sum => CSA_sum_1_27_0, c_out => CSA_carry_1_27_0);
FA_lbl_1_27_1: FA port map(in1 => CSA_sum_0_27_6, in2 => CSA_sum_0_27_5, c_in => CSA_sum_0_27_4, sum => CSA_sum_1_27_1, c_out => CSA_carry_1_27_1);
FA_lbl_1_27_2: FA port map(in1 => CSA_sum_0_27_3, in2 => CSA_sum_0_27_2, c_in => CSA_sum_0_27_1, sum => CSA_sum_1_27_2, c_out => CSA_carry_1_27_2);
FA_lbl_1_27_3: FA port map(in1 => CSA_sum_0_27_0, in2 => CSA_carry_0_26_8, c_in => CSA_carry_0_26_7, sum => CSA_sum_1_27_3, c_out => CSA_carry_1_27_3);
FA_lbl_1_27_4: FA port map(in1 => CSA_carry_0_26_6, in2 => CSA_carry_0_26_5, c_in => CSA_carry_0_26_4, sum => CSA_sum_1_27_4, c_out => CSA_carry_1_27_4);
FA_lbl_1_27_5: FA port map(in1 => CSA_carry_0_26_3, in2 => CSA_carry_0_26_2, c_in => CSA_carry_0_26_1, sum => CSA_sum_1_27_5, c_out => CSA_carry_1_27_5);
FA_lbl_1_28_0: FA port map(in1 => b_and_a(865), in2 => b_and_a(896), c_in => CSA_sum_0_28_8, sum => CSA_sum_1_28_0, c_out => CSA_carry_1_28_0);
FA_lbl_1_28_1: FA port map(in1 => CSA_sum_0_28_7, in2 => CSA_sum_0_28_6, c_in => CSA_sum_0_28_5, sum => CSA_sum_1_28_1, c_out => CSA_carry_1_28_1);
FA_lbl_1_28_2: FA port map(in1 => CSA_sum_0_28_4, in2 => CSA_sum_0_28_3, c_in => CSA_sum_0_28_2, sum => CSA_sum_1_28_2, c_out => CSA_carry_1_28_2);
FA_lbl_1_28_3: FA port map(in1 => CSA_sum_0_28_1, in2 => CSA_sum_0_28_0, c_in => CSA_carry_0_27_8, sum => CSA_sum_1_28_3, c_out => CSA_carry_1_28_3);
FA_lbl_1_28_4: FA port map(in1 => CSA_carry_0_27_7, in2 => CSA_carry_0_27_6, c_in => CSA_carry_0_27_5, sum => CSA_sum_1_28_4, c_out => CSA_carry_1_28_4);
FA_lbl_1_28_5: FA port map(in1 => CSA_carry_0_27_4, in2 => CSA_carry_0_27_3, c_in => CSA_carry_0_27_2, sum => CSA_sum_1_28_5, c_out => CSA_carry_1_28_5);
FA_lbl_1_29_0: FA port map(in1 => CSA_sum_0_29_9, in2 => CSA_sum_0_29_8, c_in => CSA_sum_0_29_7, sum => CSA_sum_1_29_0, c_out => CSA_carry_1_29_0);
FA_lbl_1_29_1: FA port map(in1 => CSA_sum_0_29_6, in2 => CSA_sum_0_29_5, c_in => CSA_sum_0_29_4, sum => CSA_sum_1_29_1, c_out => CSA_carry_1_29_1);
FA_lbl_1_29_2: FA port map(in1 => CSA_sum_0_29_3, in2 => CSA_sum_0_29_2, c_in => CSA_sum_0_29_1, sum => CSA_sum_1_29_2, c_out => CSA_carry_1_29_2);
FA_lbl_1_29_3: FA port map(in1 => CSA_sum_0_29_0, in2 => CSA_carry_0_28_8, c_in => CSA_carry_0_28_7, sum => CSA_sum_1_29_3, c_out => CSA_carry_1_29_3);
FA_lbl_1_29_4: FA port map(in1 => CSA_carry_0_28_6, in2 => CSA_carry_0_28_5, c_in => CSA_carry_0_28_4, sum => CSA_sum_1_29_4, c_out => CSA_carry_1_29_4);
FA_lbl_1_29_5: FA port map(in1 => CSA_carry_0_28_3, in2 => CSA_carry_0_28_2, c_in => CSA_carry_0_28_1, sum => CSA_sum_1_29_5, c_out => CSA_carry_1_29_5);
FA_lbl_1_30_0: FA port map(in1 => b_and_a(960), in2 => CSA_sum_0_30_9, c_in => CSA_sum_0_30_8, sum => CSA_sum_1_30_0, c_out => CSA_carry_1_30_0);
FA_lbl_1_30_1: FA port map(in1 => CSA_sum_0_30_7, in2 => CSA_sum_0_30_6, c_in => CSA_sum_0_30_5, sum => CSA_sum_1_30_1, c_out => CSA_carry_1_30_1);
FA_lbl_1_30_2: FA port map(in1 => CSA_sum_0_30_4, in2 => CSA_sum_0_30_3, c_in => CSA_sum_0_30_2, sum => CSA_sum_1_30_2, c_out => CSA_carry_1_30_2);
FA_lbl_1_30_3: FA port map(in1 => CSA_sum_0_30_1, in2 => CSA_sum_0_30_0, c_in => CSA_carry_0_29_9, sum => CSA_sum_1_30_3, c_out => CSA_carry_1_30_3);
FA_lbl_1_30_4: FA port map(in1 => CSA_carry_0_29_8, in2 => CSA_carry_0_29_7, c_in => CSA_carry_0_29_6, sum => CSA_sum_1_30_4, c_out => CSA_carry_1_30_4);
FA_lbl_1_30_5: FA port map(in1 => CSA_carry_0_29_5, in2 => CSA_carry_0_29_4, c_in => CSA_carry_0_29_3, sum => CSA_sum_1_30_5, c_out => CSA_carry_1_30_5);
FA_lbl_1_30_6: FA port map(in1 => CSA_carry_0_29_2, in2 => CSA_carry_0_29_1, c_in => CSA_carry_0_29_0, sum => CSA_sum_1_30_6, c_out => CSA_carry_1_30_6);
FA_lbl_1_31_0: FA port map(in1 => b_and_a(961), in2 => b_and_a(992), c_in => CSA_sum_0_31_9, sum => CSA_sum_1_31_0, c_out => CSA_carry_1_31_0);
FA_lbl_1_31_1: FA port map(in1 => CSA_sum_0_31_8, in2 => CSA_sum_0_31_7, c_in => CSA_sum_0_31_6, sum => CSA_sum_1_31_1, c_out => CSA_carry_1_31_1);
FA_lbl_1_31_2: FA port map(in1 => CSA_sum_0_31_5, in2 => CSA_sum_0_31_4, c_in => CSA_sum_0_31_3, sum => CSA_sum_1_31_2, c_out => CSA_carry_1_31_2);
FA_lbl_1_31_3: FA port map(in1 => CSA_sum_0_31_2, in2 => CSA_sum_0_31_1, c_in => CSA_sum_0_31_0, sum => CSA_sum_1_31_3, c_out => CSA_carry_1_31_3);
FA_lbl_1_31_4: FA port map(in1 => CSA_carry_0_30_9, in2 => CSA_carry_0_30_8, c_in => CSA_carry_0_30_7, sum => CSA_sum_1_31_4, c_out => CSA_carry_1_31_4);
FA_lbl_1_31_5: FA port map(in1 => CSA_carry_0_30_6, in2 => CSA_carry_0_30_5, c_in => CSA_carry_0_30_4, sum => CSA_sum_1_31_5, c_out => CSA_carry_1_31_5);
FA_lbl_1_31_6: FA port map(in1 => CSA_carry_0_30_3, in2 => CSA_carry_0_30_2, c_in => CSA_carry_0_30_1, sum => CSA_sum_1_31_6, c_out => CSA_carry_1_31_6);
FA_lbl_1_32_0: FA port map(in1 => b_and_a(993), in2 => CSA_sum_0_32_9, c_in => CSA_sum_0_32_8, sum => CSA_sum_1_32_0, c_out => CSA_carry_1_32_0);
FA_lbl_1_32_1: FA port map(in1 => CSA_sum_0_32_7, in2 => CSA_sum_0_32_6, c_in => CSA_sum_0_32_5, sum => CSA_sum_1_32_1, c_out => CSA_carry_1_32_1);
FA_lbl_1_32_2: FA port map(in1 => CSA_sum_0_32_4, in2 => CSA_sum_0_32_3, c_in => CSA_sum_0_32_2, sum => CSA_sum_1_32_2, c_out => CSA_carry_1_32_2);
FA_lbl_1_32_3: FA port map(in1 => CSA_sum_0_32_1, in2 => CSA_sum_0_32_0, c_in => CSA_carry_0_31_9, sum => CSA_sum_1_32_3, c_out => CSA_carry_1_32_3);
FA_lbl_1_32_4: FA port map(in1 => CSA_carry_0_31_8, in2 => CSA_carry_0_31_7, c_in => CSA_carry_0_31_6, sum => CSA_sum_1_32_4, c_out => CSA_carry_1_32_4);
FA_lbl_1_32_5: FA port map(in1 => CSA_carry_0_31_5, in2 => CSA_carry_0_31_4, c_in => CSA_carry_0_31_3, sum => CSA_sum_1_32_5, c_out => CSA_carry_1_32_5);
FA_lbl_1_32_6: FA port map(in1 => CSA_carry_0_31_2, in2 => CSA_carry_0_31_1, c_in => CSA_carry_0_31_0, sum => CSA_sum_1_32_6, c_out => CSA_carry_1_32_6);
FA_lbl_1_33_0: FA port map(in1 => CSA_sum_0_33_9, in2 => CSA_sum_0_33_8, c_in => CSA_sum_0_33_7, sum => CSA_sum_1_33_0, c_out => CSA_carry_1_33_0);
FA_lbl_1_33_1: FA port map(in1 => CSA_sum_0_33_6, in2 => CSA_sum_0_33_5, c_in => CSA_sum_0_33_4, sum => CSA_sum_1_33_1, c_out => CSA_carry_1_33_1);
FA_lbl_1_33_2: FA port map(in1 => CSA_sum_0_33_3, in2 => CSA_sum_0_33_2, c_in => CSA_sum_0_33_1, sum => CSA_sum_1_33_2, c_out => CSA_carry_1_33_2);
FA_lbl_1_33_3: FA port map(in1 => CSA_sum_0_33_0, in2 => CSA_carry_0_32_9, c_in => CSA_carry_0_32_8, sum => CSA_sum_1_33_3, c_out => CSA_carry_1_33_3);
FA_lbl_1_33_4: FA port map(in1 => CSA_carry_0_32_7, in2 => CSA_carry_0_32_6, c_in => CSA_carry_0_32_5, sum => CSA_sum_1_33_4, c_out => CSA_carry_1_33_4);
FA_lbl_1_33_5: FA port map(in1 => CSA_carry_0_32_4, in2 => CSA_carry_0_32_3, c_in => CSA_carry_0_32_2, sum => CSA_sum_1_33_5, c_out => CSA_carry_1_33_5);
FA_lbl_1_34_0: FA port map(in1 => b_and_a(964), in2 => b_and_a(995), c_in => CSA_sum_0_34_8, sum => CSA_sum_1_34_0, c_out => CSA_carry_1_34_0);
FA_lbl_1_34_1: FA port map(in1 => CSA_sum_0_34_7, in2 => CSA_sum_0_34_6, c_in => CSA_sum_0_34_5, sum => CSA_sum_1_34_1, c_out => CSA_carry_1_34_1);
FA_lbl_1_34_2: FA port map(in1 => CSA_sum_0_34_4, in2 => CSA_sum_0_34_3, c_in => CSA_sum_0_34_2, sum => CSA_sum_1_34_2, c_out => CSA_carry_1_34_2);
FA_lbl_1_34_3: FA port map(in1 => CSA_sum_0_34_1, in2 => CSA_sum_0_34_0, c_in => CSA_carry_0_33_9, sum => CSA_sum_1_34_3, c_out => CSA_carry_1_34_3);
FA_lbl_1_34_4: FA port map(in1 => CSA_carry_0_33_8, in2 => CSA_carry_0_33_7, c_in => CSA_carry_0_33_6, sum => CSA_sum_1_34_4, c_out => CSA_carry_1_34_4);
FA_lbl_1_34_5: FA port map(in1 => CSA_carry_0_33_5, in2 => CSA_carry_0_33_4, c_in => CSA_carry_0_33_3, sum => CSA_sum_1_34_5, c_out => CSA_carry_1_34_5);
FA_lbl_1_34_6: FA port map(in1 => CSA_carry_0_33_2, in2 => CSA_carry_0_33_1, c_in => CSA_carry_0_33_0, sum => CSA_sum_1_34_6, c_out => CSA_carry_1_34_6);
FA_lbl_1_35_0: FA port map(in1 => b_and_a(996), in2 => CSA_sum_0_35_8, c_in => CSA_sum_0_35_7, sum => CSA_sum_1_35_0, c_out => CSA_carry_1_35_0);
FA_lbl_1_35_1: FA port map(in1 => CSA_sum_0_35_6, in2 => CSA_sum_0_35_5, c_in => CSA_sum_0_35_4, sum => CSA_sum_1_35_1, c_out => CSA_carry_1_35_1);
FA_lbl_1_35_2: FA port map(in1 => CSA_sum_0_35_3, in2 => CSA_sum_0_35_2, c_in => CSA_sum_0_35_1, sum => CSA_sum_1_35_2, c_out => CSA_carry_1_35_2);
FA_lbl_1_35_3: FA port map(in1 => CSA_sum_0_35_0, in2 => CSA_carry_0_34_8, c_in => CSA_carry_0_34_7, sum => CSA_sum_1_35_3, c_out => CSA_carry_1_35_3);
FA_lbl_1_35_4: FA port map(in1 => CSA_carry_0_34_6, in2 => CSA_carry_0_34_5, c_in => CSA_carry_0_34_4, sum => CSA_sum_1_35_4, c_out => CSA_carry_1_35_4);
FA_lbl_1_35_5: FA port map(in1 => CSA_carry_0_34_3, in2 => CSA_carry_0_34_2, c_in => CSA_carry_0_34_1, sum => CSA_sum_1_35_5, c_out => CSA_carry_1_35_5);
FA_lbl_1_36_0: FA port map(in1 => CSA_sum_0_36_8, in2 => CSA_sum_0_36_7, c_in => CSA_sum_0_36_6, sum => CSA_sum_1_36_0, c_out => CSA_carry_1_36_0);
FA_lbl_1_36_1: FA port map(in1 => CSA_sum_0_36_5, in2 => CSA_sum_0_36_4, c_in => CSA_sum_0_36_3, sum => CSA_sum_1_36_1, c_out => CSA_carry_1_36_1);
FA_lbl_1_36_2: FA port map(in1 => CSA_sum_0_36_2, in2 => CSA_sum_0_36_1, c_in => CSA_sum_0_36_0, sum => CSA_sum_1_36_2, c_out => CSA_carry_1_36_2);
FA_lbl_1_36_3: FA port map(in1 => CSA_carry_0_35_8, in2 => CSA_carry_0_35_7, c_in => CSA_carry_0_35_6, sum => CSA_sum_1_36_3, c_out => CSA_carry_1_36_3);
FA_lbl_1_36_4: FA port map(in1 => CSA_carry_0_35_5, in2 => CSA_carry_0_35_4, c_in => CSA_carry_0_35_3, sum => CSA_sum_1_36_4, c_out => CSA_carry_1_36_4);
FA_lbl_1_36_5: FA port map(in1 => CSA_carry_0_35_2, in2 => CSA_carry_0_35_1, c_in => CSA_carry_0_35_0, sum => CSA_sum_1_36_5, c_out => CSA_carry_1_36_5);
FA_lbl_1_37_0: FA port map(in1 => b_and_a(967), in2 => b_and_a(998), c_in => CSA_sum_0_37_7, sum => CSA_sum_1_37_0, c_out => CSA_carry_1_37_0);
FA_lbl_1_37_1: FA port map(in1 => CSA_sum_0_37_6, in2 => CSA_sum_0_37_5, c_in => CSA_sum_0_37_4, sum => CSA_sum_1_37_1, c_out => CSA_carry_1_37_1);
FA_lbl_1_37_2: FA port map(in1 => CSA_sum_0_37_3, in2 => CSA_sum_0_37_2, c_in => CSA_sum_0_37_1, sum => CSA_sum_1_37_2, c_out => CSA_carry_1_37_2);
FA_lbl_1_37_3: FA port map(in1 => CSA_sum_0_37_0, in2 => CSA_carry_0_36_8, c_in => CSA_carry_0_36_7, sum => CSA_sum_1_37_3, c_out => CSA_carry_1_37_3);
FA_lbl_1_37_4: FA port map(in1 => CSA_carry_0_36_6, in2 => CSA_carry_0_36_5, c_in => CSA_carry_0_36_4, sum => CSA_sum_1_37_4, c_out => CSA_carry_1_37_4);
FA_lbl_1_37_5: FA port map(in1 => CSA_carry_0_36_3, in2 => CSA_carry_0_36_2, c_in => CSA_carry_0_36_1, sum => CSA_sum_1_37_5, c_out => CSA_carry_1_37_5);
FA_lbl_1_38_0: FA port map(in1 => b_and_a(999), in2 => CSA_sum_0_38_7, c_in => CSA_sum_0_38_6, sum => CSA_sum_1_38_0, c_out => CSA_carry_1_38_0);
FA_lbl_1_38_1: FA port map(in1 => CSA_sum_0_38_5, in2 => CSA_sum_0_38_4, c_in => CSA_sum_0_38_3, sum => CSA_sum_1_38_1, c_out => CSA_carry_1_38_1);
FA_lbl_1_38_2: FA port map(in1 => CSA_sum_0_38_2, in2 => CSA_sum_0_38_1, c_in => CSA_sum_0_38_0, sum => CSA_sum_1_38_2, c_out => CSA_carry_1_38_2);
FA_lbl_1_38_3: FA port map(in1 => CSA_carry_0_37_7, in2 => CSA_carry_0_37_6, c_in => CSA_carry_0_37_5, sum => CSA_sum_1_38_3, c_out => CSA_carry_1_38_3);
FA_lbl_1_38_4: FA port map(in1 => CSA_carry_0_37_4, in2 => CSA_carry_0_37_3, c_in => CSA_carry_0_37_2, sum => CSA_sum_1_38_4, c_out => CSA_carry_1_38_4);
FA_lbl_1_39_0: FA port map(in1 => CSA_sum_0_39_7, in2 => CSA_sum_0_39_6, c_in => CSA_sum_0_39_5, sum => CSA_sum_1_39_0, c_out => CSA_carry_1_39_0);
FA_lbl_1_39_1: FA port map(in1 => CSA_sum_0_39_4, in2 => CSA_sum_0_39_3, c_in => CSA_sum_0_39_2, sum => CSA_sum_1_39_1, c_out => CSA_carry_1_39_1);
FA_lbl_1_39_2: FA port map(in1 => CSA_sum_0_39_1, in2 => CSA_sum_0_39_0, c_in => CSA_carry_0_38_7, sum => CSA_sum_1_39_2, c_out => CSA_carry_1_39_2);
FA_lbl_1_39_3: FA port map(in1 => CSA_carry_0_38_6, in2 => CSA_carry_0_38_5, c_in => CSA_carry_0_38_4, sum => CSA_sum_1_39_3, c_out => CSA_carry_1_39_3);
FA_lbl_1_39_4: FA port map(in1 => CSA_carry_0_38_3, in2 => CSA_carry_0_38_2, c_in => CSA_carry_0_38_1, sum => CSA_sum_1_39_4, c_out => CSA_carry_1_39_4);
FA_lbl_1_40_0: FA port map(in1 => b_and_a(970), in2 => b_and_a(1001), c_in => CSA_sum_0_40_6, sum => CSA_sum_1_40_0, c_out => CSA_carry_1_40_0);
FA_lbl_1_40_1: FA port map(in1 => CSA_sum_0_40_5, in2 => CSA_sum_0_40_4, c_in => CSA_sum_0_40_3, sum => CSA_sum_1_40_1, c_out => CSA_carry_1_40_1);
FA_lbl_1_40_2: FA port map(in1 => CSA_sum_0_40_2, in2 => CSA_sum_0_40_1, c_in => CSA_sum_0_40_0, sum => CSA_sum_1_40_2, c_out => CSA_carry_1_40_2);
FA_lbl_1_40_3: FA port map(in1 => CSA_carry_0_39_7, in2 => CSA_carry_0_39_6, c_in => CSA_carry_0_39_5, sum => CSA_sum_1_40_3, c_out => CSA_carry_1_40_3);
FA_lbl_1_40_4: FA port map(in1 => CSA_carry_0_39_4, in2 => CSA_carry_0_39_3, c_in => CSA_carry_0_39_2, sum => CSA_sum_1_40_4, c_out => CSA_carry_1_40_4);
FA_lbl_1_41_0: FA port map(in1 => b_and_a(1002), in2 => CSA_sum_0_41_6, c_in => CSA_sum_0_41_5, sum => CSA_sum_1_41_0, c_out => CSA_carry_1_41_0);
FA_lbl_1_41_1: FA port map(in1 => CSA_sum_0_41_4, in2 => CSA_sum_0_41_3, c_in => CSA_sum_0_41_2, sum => CSA_sum_1_41_1, c_out => CSA_carry_1_41_1);
FA_lbl_1_41_2: FA port map(in1 => CSA_sum_0_41_1, in2 => CSA_sum_0_41_0, c_in => CSA_carry_0_40_6, sum => CSA_sum_1_41_2, c_out => CSA_carry_1_41_2);
FA_lbl_1_41_3: FA port map(in1 => CSA_carry_0_40_5, in2 => CSA_carry_0_40_4, c_in => CSA_carry_0_40_3, sum => CSA_sum_1_41_3, c_out => CSA_carry_1_41_3);
FA_lbl_1_41_4: FA port map(in1 => CSA_carry_0_40_2, in2 => CSA_carry_0_40_1, c_in => CSA_carry_0_40_0, sum => CSA_sum_1_41_4, c_out => CSA_carry_1_41_4);
FA_lbl_1_42_0: FA port map(in1 => CSA_sum_0_42_6, in2 => CSA_sum_0_42_5, c_in => CSA_sum_0_42_4, sum => CSA_sum_1_42_0, c_out => CSA_carry_1_42_0);
FA_lbl_1_42_1: FA port map(in1 => CSA_sum_0_42_3, in2 => CSA_sum_0_42_2, c_in => CSA_sum_0_42_1, sum => CSA_sum_1_42_1, c_out => CSA_carry_1_42_1);
FA_lbl_1_42_2: FA port map(in1 => CSA_sum_0_42_0, in2 => CSA_carry_0_41_6, c_in => CSA_carry_0_41_5, sum => CSA_sum_1_42_2, c_out => CSA_carry_1_42_2);
FA_lbl_1_42_3: FA port map(in1 => CSA_carry_0_41_4, in2 => CSA_carry_0_41_3, c_in => CSA_carry_0_41_2, sum => CSA_sum_1_42_3, c_out => CSA_carry_1_42_3);
FA_lbl_1_43_0: FA port map(in1 => b_and_a(973), in2 => b_and_a(1004), c_in => CSA_sum_0_43_5, sum => CSA_sum_1_43_0, c_out => CSA_carry_1_43_0);
FA_lbl_1_43_1: FA port map(in1 => CSA_sum_0_43_4, in2 => CSA_sum_0_43_3, c_in => CSA_sum_0_43_2, sum => CSA_sum_1_43_1, c_out => CSA_carry_1_43_1);
FA_lbl_1_43_2: FA port map(in1 => CSA_sum_0_43_1, in2 => CSA_sum_0_43_0, c_in => CSA_carry_0_42_6, sum => CSA_sum_1_43_2, c_out => CSA_carry_1_43_2);
FA_lbl_1_43_3: FA port map(in1 => CSA_carry_0_42_5, in2 => CSA_carry_0_42_4, c_in => CSA_carry_0_42_3, sum => CSA_sum_1_43_3, c_out => CSA_carry_1_43_3);
FA_lbl_1_43_4: FA port map(in1 => CSA_carry_0_42_2, in2 => CSA_carry_0_42_1, c_in => CSA_carry_0_42_0, sum => CSA_sum_1_43_4, c_out => CSA_carry_1_43_4);
FA_lbl_1_44_0: FA port map(in1 => b_and_a(1005), in2 => CSA_sum_0_44_5, c_in => CSA_sum_0_44_4, sum => CSA_sum_1_44_0, c_out => CSA_carry_1_44_0);
FA_lbl_1_44_1: FA port map(in1 => CSA_sum_0_44_3, in2 => CSA_sum_0_44_2, c_in => CSA_sum_0_44_1, sum => CSA_sum_1_44_1, c_out => CSA_carry_1_44_1);
FA_lbl_1_44_2: FA port map(in1 => CSA_sum_0_44_0, in2 => CSA_carry_0_43_5, c_in => CSA_carry_0_43_4, sum => CSA_sum_1_44_2, c_out => CSA_carry_1_44_2);
FA_lbl_1_44_3: FA port map(in1 => CSA_carry_0_43_3, in2 => CSA_carry_0_43_2, c_in => CSA_carry_0_43_1, sum => CSA_sum_1_44_3, c_out => CSA_carry_1_44_3);
FA_lbl_1_45_0: FA port map(in1 => CSA_sum_0_45_5, in2 => CSA_sum_0_45_4, c_in => CSA_sum_0_45_3, sum => CSA_sum_1_45_0, c_out => CSA_carry_1_45_0);
FA_lbl_1_45_1: FA port map(in1 => CSA_sum_0_45_2, in2 => CSA_sum_0_45_1, c_in => CSA_sum_0_45_0, sum => CSA_sum_1_45_1, c_out => CSA_carry_1_45_1);
FA_lbl_1_45_2: FA port map(in1 => CSA_carry_0_44_5, in2 => CSA_carry_0_44_4, c_in => CSA_carry_0_44_3, sum => CSA_sum_1_45_2, c_out => CSA_carry_1_45_2);
FA_lbl_1_45_3: FA port map(in1 => CSA_carry_0_44_2, in2 => CSA_carry_0_44_1, c_in => CSA_carry_0_44_0, sum => CSA_sum_1_45_3, c_out => CSA_carry_1_45_3);
FA_lbl_1_46_0: FA port map(in1 => b_and_a(976), in2 => b_and_a(1007), c_in => CSA_sum_0_46_4, sum => CSA_sum_1_46_0, c_out => CSA_carry_1_46_0);
FA_lbl_1_46_1: FA port map(in1 => CSA_sum_0_46_3, in2 => CSA_sum_0_46_2, c_in => CSA_sum_0_46_1, sum => CSA_sum_1_46_1, c_out => CSA_carry_1_46_1);
FA_lbl_1_46_2: FA port map(in1 => CSA_sum_0_46_0, in2 => CSA_carry_0_45_5, c_in => CSA_carry_0_45_4, sum => CSA_sum_1_46_2, c_out => CSA_carry_1_46_2);
FA_lbl_1_46_3: FA port map(in1 => CSA_carry_0_45_3, in2 => CSA_carry_0_45_2, c_in => CSA_carry_0_45_1, sum => CSA_sum_1_46_3, c_out => CSA_carry_1_46_3);
FA_lbl_1_47_0: FA port map(in1 => b_and_a(1008), in2 => CSA_sum_0_47_4, c_in => CSA_sum_0_47_3, sum => CSA_sum_1_47_0, c_out => CSA_carry_1_47_0);
FA_lbl_1_47_1: FA port map(in1 => CSA_sum_0_47_2, in2 => CSA_sum_0_47_1, c_in => CSA_sum_0_47_0, sum => CSA_sum_1_47_1, c_out => CSA_carry_1_47_1);
FA_lbl_1_47_2: FA port map(in1 => CSA_carry_0_46_4, in2 => CSA_carry_0_46_3, c_in => CSA_carry_0_46_2, sum => CSA_sum_1_47_2, c_out => CSA_carry_1_47_2);
FA_lbl_1_48_0: FA port map(in1 => CSA_sum_0_48_4, in2 => CSA_sum_0_48_3, c_in => CSA_sum_0_48_2, sum => CSA_sum_1_48_0, c_out => CSA_carry_1_48_0);
FA_lbl_1_48_1: FA port map(in1 => CSA_sum_0_48_1, in2 => CSA_sum_0_48_0, c_in => CSA_carry_0_47_4, sum => CSA_sum_1_48_1, c_out => CSA_carry_1_48_1);
FA_lbl_1_48_2: FA port map(in1 => CSA_carry_0_47_3, in2 => CSA_carry_0_47_2, c_in => CSA_carry_0_47_1, sum => CSA_sum_1_48_2, c_out => CSA_carry_1_48_2);
FA_lbl_1_49_0: FA port map(in1 => b_and_a(979), in2 => b_and_a(1010), c_in => CSA_sum_0_49_3, sum => CSA_sum_1_49_0, c_out => CSA_carry_1_49_0);
FA_lbl_1_49_1: FA port map(in1 => CSA_sum_0_49_2, in2 => CSA_sum_0_49_1, c_in => CSA_sum_0_49_0, sum => CSA_sum_1_49_1, c_out => CSA_carry_1_49_1);
FA_lbl_1_49_2: FA port map(in1 => CSA_carry_0_48_4, in2 => CSA_carry_0_48_3, c_in => CSA_carry_0_48_2, sum => CSA_sum_1_49_2, c_out => CSA_carry_1_49_2);
FA_lbl_1_50_0: FA port map(in1 => b_and_a(1011), in2 => CSA_sum_0_50_3, c_in => CSA_sum_0_50_2, sum => CSA_sum_1_50_0, c_out => CSA_carry_1_50_0);
FA_lbl_1_50_1: FA port map(in1 => CSA_sum_0_50_1, in2 => CSA_sum_0_50_0, c_in => CSA_carry_0_49_3, sum => CSA_sum_1_50_1, c_out => CSA_carry_1_50_1);
FA_lbl_1_50_2: FA port map(in1 => CSA_carry_0_49_2, in2 => CSA_carry_0_49_1, c_in => CSA_carry_0_49_0, sum => CSA_sum_1_50_2, c_out => CSA_carry_1_50_2);
FA_lbl_1_51_0: FA port map(in1 => CSA_sum_0_51_3, in2 => CSA_sum_0_51_2, c_in => CSA_sum_0_51_1, sum => CSA_sum_1_51_0, c_out => CSA_carry_1_51_0);
FA_lbl_1_51_1: FA port map(in1 => CSA_sum_0_51_0, in2 => CSA_carry_0_50_3, c_in => CSA_carry_0_50_2, sum => CSA_sum_1_51_1, c_out => CSA_carry_1_51_1);
FA_lbl_1_52_0: FA port map(in1 => b_and_a(982), in2 => b_and_a(1013), c_in => CSA_sum_0_52_2, sum => CSA_sum_1_52_0, c_out => CSA_carry_1_52_0);
FA_lbl_1_52_1: FA port map(in1 => CSA_sum_0_52_1, in2 => CSA_sum_0_52_0, c_in => CSA_carry_0_51_3, sum => CSA_sum_1_52_1, c_out => CSA_carry_1_52_1);
FA_lbl_1_52_2: FA port map(in1 => CSA_carry_0_51_2, in2 => CSA_carry_0_51_1, c_in => CSA_carry_0_51_0, sum => CSA_sum_1_52_2, c_out => CSA_carry_1_52_2);
FA_lbl_1_53_0: FA port map(in1 => b_and_a(1014), in2 => CSA_sum_0_53_2, c_in => CSA_sum_0_53_1, sum => CSA_sum_1_53_0, c_out => CSA_carry_1_53_0);
FA_lbl_1_53_1: FA port map(in1 => CSA_sum_0_53_0, in2 => CSA_carry_0_52_2, c_in => CSA_carry_0_52_1, sum => CSA_sum_1_53_1, c_out => CSA_carry_1_53_1);
FA_lbl_1_54_0: FA port map(in1 => CSA_sum_0_54_2, in2 => CSA_sum_0_54_1, c_in => CSA_sum_0_54_0, sum => CSA_sum_1_54_0, c_out => CSA_carry_1_54_0);
FA_lbl_1_54_1: FA port map(in1 => CSA_carry_0_53_2, in2 => CSA_carry_0_53_1, c_in => CSA_carry_0_53_0, sum => CSA_sum_1_54_1, c_out => CSA_carry_1_54_1);
FA_lbl_1_55_0: FA port map(in1 => b_and_a(985), in2 => b_and_a(1016), c_in => CSA_sum_0_55_1, sum => CSA_sum_1_55_0, c_out => CSA_carry_1_55_0);
FA_lbl_1_55_1: FA port map(in1 => CSA_sum_0_55_0, in2 => CSA_carry_0_54_2, c_in => CSA_carry_0_54_1, sum => CSA_sum_1_55_1, c_out => CSA_carry_1_55_1);
FA_lbl_1_56_0: FA port map(in1 => b_and_a(1017), in2 => CSA_sum_0_56_1, c_in => CSA_sum_0_56_0, sum => CSA_sum_1_56_0, c_out => CSA_carry_1_56_0);
FA_lbl_1_57_0: FA port map(in1 => CSA_sum_0_57_1, in2 => CSA_sum_0_57_0, c_in => CSA_carry_0_56_1, sum => CSA_sum_1_57_0, c_out => CSA_carry_1_57_0);
FA_lbl_1_58_0: FA port map(in1 => b_and_a(988), in2 => b_and_a(1019), c_in => CSA_sum_0_58_0, sum => CSA_sum_1_58_0, c_out => CSA_carry_1_58_0);
FA_lbl_1_59_0: FA port map(in1 => b_and_a(1020), in2 => CSA_sum_0_59_0, c_in => CSA_carry_0_58_0, sum => CSA_sum_1_59_0, c_out => CSA_carry_1_59_0);
FA_lbl_1_61_0: FA port map(in1 => b_and_a(991), in2 => b_and_a(1022), c_in => CSA_carry_0_60_0, sum => CSA_sum_1_61_0, c_out => CSA_carry_1_61_0);
FA_lbl_2_4_0: FA port map(in1 => CSA_sum_1_4_0, in2 => CSA_carry_1_3_0, c_in => CSA_carry_0_3_0, sum => CSA_sum_2_4_0, c_out => CSA_carry_2_4_0);
FA_lbl_2_6_0: FA port map(in1 => CSA_sum_1_6_0, in2 => CSA_carry_1_5_0, c_in => CSA_carry_0_5_1, sum => CSA_sum_2_6_0, c_out => CSA_carry_2_6_0);
FA_lbl_2_7_0: FA port map(in1 => CSA_sum_1_7_1, in2 => CSA_sum_1_7_0, c_in => CSA_carry_1_6_0, sum => CSA_sum_2_7_0, c_out => CSA_carry_2_7_0);
FA_lbl_2_8_0: FA port map(in1 => CSA_sum_1_8_0, in2 => CSA_carry_1_7_1, c_in => CSA_carry_1_7_0, sum => CSA_sum_2_8_0, c_out => CSA_carry_2_8_0);
FA_lbl_2_9_0: FA port map(in1 => CSA_sum_1_9_1, in2 => CSA_sum_1_9_0, c_in => CSA_carry_1_8_0, sum => CSA_sum_2_9_0, c_out => CSA_carry_2_9_0);
FA_lbl_2_10_0: FA port map(in1 => CSA_sum_1_10_1, in2 => CSA_sum_1_10_0, c_in => CSA_carry_1_9_1, sum => CSA_sum_2_10_0, c_out => CSA_carry_2_10_0);
FA_lbl_2_10_1: FA port map(in1 => CSA_carry_1_9_0, in2 => CSA_carry_0_9_1, c_in => CSA_carry_0_9_0, sum => CSA_sum_2_10_1, c_out => CSA_carry_2_10_1);
FA_lbl_2_11_0: FA port map(in1 => CSA_sum_1_11_1, in2 => CSA_sum_1_11_0, c_in => CSA_carry_1_10_1, sum => CSA_sum_2_11_0, c_out => CSA_carry_2_11_0);
FA_lbl_2_12_0: FA port map(in1 => CSA_sum_1_12_2, in2 => CSA_sum_1_12_1, c_in => CSA_sum_1_12_0, sum => CSA_sum_2_12_0, c_out => CSA_carry_2_12_0);
FA_lbl_2_13_0: FA port map(in1 => CSA_sum_1_13_2, in2 => CSA_sum_1_13_1, c_in => CSA_sum_1_13_0, sum => CSA_sum_2_13_0, c_out => CSA_carry_2_13_0);
FA_lbl_2_13_1: FA port map(in1 => CSA_carry_1_12_2, in2 => CSA_carry_1_12_1, c_in => CSA_carry_1_12_0, sum => CSA_sum_2_13_1, c_out => CSA_carry_2_13_1);
FA_lbl_2_14_0: FA port map(in1 => CSA_sum_1_14_2, in2 => CSA_sum_1_14_1, c_in => CSA_sum_1_14_0, sum => CSA_sum_2_14_0, c_out => CSA_carry_2_14_0);
FA_lbl_2_14_1: FA port map(in1 => CSA_carry_1_13_2, in2 => CSA_carry_1_13_1, c_in => CSA_carry_1_13_0, sum => CSA_sum_2_14_1, c_out => CSA_carry_2_14_1);
FA_lbl_2_15_0: FA port map(in1 => CSA_sum_1_15_2, in2 => CSA_sum_1_15_1, c_in => CSA_sum_1_15_0, sum => CSA_sum_2_15_0, c_out => CSA_carry_2_15_0);
FA_lbl_2_15_1: FA port map(in1 => CSA_carry_1_14_2, in2 => CSA_carry_1_14_1, c_in => CSA_carry_1_14_0, sum => CSA_sum_2_15_1, c_out => CSA_carry_2_15_1);
FA_lbl_2_16_0: FA port map(in1 => CSA_sum_1_16_3, in2 => CSA_sum_1_16_2, c_in => CSA_sum_1_16_1, sum => CSA_sum_2_16_0, c_out => CSA_carry_2_16_0);
FA_lbl_2_16_1: FA port map(in1 => CSA_sum_1_16_0, in2 => CSA_carry_1_15_2, c_in => CSA_carry_1_15_1, sum => CSA_sum_2_16_1, c_out => CSA_carry_2_16_1);
FA_lbl_2_17_0: FA port map(in1 => CSA_sum_1_17_2, in2 => CSA_sum_1_17_1, c_in => CSA_sum_1_17_0, sum => CSA_sum_2_17_0, c_out => CSA_carry_2_17_0);
FA_lbl_2_17_1: FA port map(in1 => CSA_carry_1_16_3, in2 => CSA_carry_1_16_2, c_in => CSA_carry_1_16_1, sum => CSA_sum_2_17_1, c_out => CSA_carry_2_17_1);
FA_lbl_2_17_2: FA port map(in1 => CSA_carry_1_16_0, in2 => CSA_carry_0_16_1, c_in => CSA_carry_0_16_0, sum => CSA_sum_2_17_2, c_out => CSA_carry_2_17_2);
FA_lbl_2_18_0: FA port map(in1 => CSA_sum_1_18_3, in2 => CSA_sum_1_18_2, c_in => CSA_sum_1_18_1, sum => CSA_sum_2_18_0, c_out => CSA_carry_2_18_0);
FA_lbl_2_18_1: FA port map(in1 => CSA_sum_1_18_0, in2 => CSA_carry_1_17_2, c_in => CSA_carry_1_17_1, sum => CSA_sum_2_18_1, c_out => CSA_carry_2_18_1);
FA_lbl_2_19_0: FA port map(in1 => CSA_sum_1_19_3, in2 => CSA_sum_1_19_2, c_in => CSA_sum_1_19_1, sum => CSA_sum_2_19_0, c_out => CSA_carry_2_19_0);
FA_lbl_2_19_1: FA port map(in1 => CSA_sum_1_19_0, in2 => CSA_carry_1_18_3, c_in => CSA_carry_1_18_2, sum => CSA_sum_2_19_1, c_out => CSA_carry_2_19_1);
FA_lbl_2_19_2: FA port map(in1 => CSA_carry_1_18_1, in2 => CSA_carry_1_18_0, c_in => CSA_carry_0_18_1, sum => CSA_sum_2_19_2, c_out => CSA_carry_2_19_2);
FA_lbl_2_20_0: FA port map(in1 => CSA_sum_1_20_3, in2 => CSA_sum_1_20_2, c_in => CSA_sum_1_20_1, sum => CSA_sum_2_20_0, c_out => CSA_carry_2_20_0);
FA_lbl_2_20_1: FA port map(in1 => CSA_sum_1_20_0, in2 => CSA_carry_1_19_3, c_in => CSA_carry_1_19_2, sum => CSA_sum_2_20_1, c_out => CSA_carry_2_20_1);
FA_lbl_2_20_2: FA port map(in1 => CSA_carry_1_19_1, in2 => CSA_carry_1_19_0, c_in => CSA_carry_0_19_0, sum => CSA_sum_2_20_2, c_out => CSA_carry_2_20_2);
FA_lbl_2_21_0: FA port map(in1 => CSA_sum_1_21_4, in2 => CSA_sum_1_21_3, c_in => CSA_sum_1_21_2, sum => CSA_sum_2_21_0, c_out => CSA_carry_2_21_0);
FA_lbl_2_21_1: FA port map(in1 => CSA_sum_1_21_1, in2 => CSA_sum_1_21_0, c_in => CSA_carry_1_20_3, sum => CSA_sum_2_21_1, c_out => CSA_carry_2_21_1);
FA_lbl_2_21_2: FA port map(in1 => CSA_carry_1_20_2, in2 => CSA_carry_1_20_1, c_in => CSA_carry_1_20_0, sum => CSA_sum_2_21_2, c_out => CSA_carry_2_21_2);
FA_lbl_2_22_0: FA port map(in1 => CSA_sum_1_22_4, in2 => CSA_sum_1_22_3, c_in => CSA_sum_1_22_2, sum => CSA_sum_2_22_0, c_out => CSA_carry_2_22_0);
FA_lbl_2_22_1: FA port map(in1 => CSA_sum_1_22_1, in2 => CSA_sum_1_22_0, c_in => CSA_carry_1_21_4, sum => CSA_sum_2_22_1, c_out => CSA_carry_2_22_1);
FA_lbl_2_22_2: FA port map(in1 => CSA_carry_1_21_3, in2 => CSA_carry_1_21_2, c_in => CSA_carry_1_21_1, sum => CSA_sum_2_22_2, c_out => CSA_carry_2_22_2);
FA_lbl_2_23_0: FA port map(in1 => CSA_sum_1_23_4, in2 => CSA_sum_1_23_3, c_in => CSA_sum_1_23_2, sum => CSA_sum_2_23_0, c_out => CSA_carry_2_23_0);
FA_lbl_2_23_1: FA port map(in1 => CSA_sum_1_23_1, in2 => CSA_sum_1_23_0, c_in => CSA_carry_1_22_4, sum => CSA_sum_2_23_1, c_out => CSA_carry_2_23_1);
FA_lbl_2_23_2: FA port map(in1 => CSA_carry_1_22_3, in2 => CSA_carry_1_22_2, c_in => CSA_carry_1_22_1, sum => CSA_sum_2_23_2, c_out => CSA_carry_2_23_2);
FA_lbl_2_24_0: FA port map(in1 => CSA_sum_1_24_4, in2 => CSA_sum_1_24_3, c_in => CSA_sum_1_24_2, sum => CSA_sum_2_24_0, c_out => CSA_carry_2_24_0);
FA_lbl_2_24_1: FA port map(in1 => CSA_sum_1_24_1, in2 => CSA_sum_1_24_0, c_in => CSA_carry_1_23_4, sum => CSA_sum_2_24_1, c_out => CSA_carry_2_24_1);
FA_lbl_2_24_2: FA port map(in1 => CSA_carry_1_23_3, in2 => CSA_carry_1_23_2, c_in => CSA_carry_1_23_1, sum => CSA_sum_2_24_2, c_out => CSA_carry_2_24_2);
FA_lbl_2_24_3: FA port map(in1 => CSA_carry_1_23_0, in2 => CSA_carry_0_23_1, c_in => CSA_carry_0_23_0, sum => CSA_sum_2_24_3, c_out => CSA_carry_2_24_3);
FA_lbl_2_25_0: FA port map(in1 => CSA_sum_1_25_5, in2 => CSA_sum_1_25_4, c_in => CSA_sum_1_25_3, sum => CSA_sum_2_25_0, c_out => CSA_carry_2_25_0);
FA_lbl_2_25_1: FA port map(in1 => CSA_sum_1_25_2, in2 => CSA_sum_1_25_1, c_in => CSA_sum_1_25_0, sum => CSA_sum_2_25_1, c_out => CSA_carry_2_25_1);
FA_lbl_2_25_2: FA port map(in1 => CSA_carry_1_24_4, in2 => CSA_carry_1_24_3, c_in => CSA_carry_1_24_2, sum => CSA_sum_2_25_2, c_out => CSA_carry_2_25_2);
FA_lbl_2_26_0: FA port map(in1 => CSA_sum_1_26_4, in2 => CSA_sum_1_26_3, c_in => CSA_sum_1_26_2, sum => CSA_sum_2_26_0, c_out => CSA_carry_2_26_0);
FA_lbl_2_26_1: FA port map(in1 => CSA_sum_1_26_1, in2 => CSA_sum_1_26_0, c_in => CSA_carry_1_25_5, sum => CSA_sum_2_26_1, c_out => CSA_carry_2_26_1);
FA_lbl_2_26_2: FA port map(in1 => CSA_carry_1_25_4, in2 => CSA_carry_1_25_3, c_in => CSA_carry_1_25_2, sum => CSA_sum_2_26_2, c_out => CSA_carry_2_26_2);
FA_lbl_2_26_3: FA port map(in1 => CSA_carry_1_25_1, in2 => CSA_carry_1_25_0, c_in => CSA_carry_0_25_1, sum => CSA_sum_2_26_3, c_out => CSA_carry_2_26_3);
FA_lbl_2_27_0: FA port map(in1 => CSA_sum_1_27_5, in2 => CSA_sum_1_27_4, c_in => CSA_sum_1_27_3, sum => CSA_sum_2_27_0, c_out => CSA_carry_2_27_0);
FA_lbl_2_27_1: FA port map(in1 => CSA_sum_1_27_2, in2 => CSA_sum_1_27_1, c_in => CSA_sum_1_27_0, sum => CSA_sum_2_27_1, c_out => CSA_carry_2_27_1);
FA_lbl_2_27_2: FA port map(in1 => CSA_carry_1_26_4, in2 => CSA_carry_1_26_3, c_in => CSA_carry_1_26_2, sum => CSA_sum_2_27_2, c_out => CSA_carry_2_27_2);
FA_lbl_2_27_3: FA port map(in1 => CSA_carry_1_26_1, in2 => CSA_carry_1_26_0, c_in => CSA_carry_0_26_0, sum => CSA_sum_2_27_3, c_out => CSA_carry_2_27_3);
FA_lbl_2_28_0: FA port map(in1 => CSA_sum_1_28_5, in2 => CSA_sum_1_28_4, c_in => CSA_sum_1_28_3, sum => CSA_sum_2_28_0, c_out => CSA_carry_2_28_0);
FA_lbl_2_28_1: FA port map(in1 => CSA_sum_1_28_2, in2 => CSA_sum_1_28_1, c_in => CSA_sum_1_28_0, sum => CSA_sum_2_28_1, c_out => CSA_carry_2_28_1);
FA_lbl_2_28_2: FA port map(in1 => CSA_carry_1_27_5, in2 => CSA_carry_1_27_4, c_in => CSA_carry_1_27_3, sum => CSA_sum_2_28_2, c_out => CSA_carry_2_28_2);
FA_lbl_2_28_3: FA port map(in1 => CSA_carry_1_27_2, in2 => CSA_carry_1_27_1, c_in => CSA_carry_1_27_0, sum => CSA_sum_2_28_3, c_out => CSA_carry_2_28_3);
FA_lbl_2_29_0: FA port map(in1 => CSA_sum_1_29_5, in2 => CSA_sum_1_29_4, c_in => CSA_sum_1_29_3, sum => CSA_sum_2_29_0, c_out => CSA_carry_2_29_0);
FA_lbl_2_29_1: FA port map(in1 => CSA_sum_1_29_2, in2 => CSA_sum_1_29_1, c_in => CSA_sum_1_29_0, sum => CSA_sum_2_29_1, c_out => CSA_carry_2_29_1);
FA_lbl_2_29_2: FA port map(in1 => CSA_carry_1_28_5, in2 => CSA_carry_1_28_4, c_in => CSA_carry_1_28_3, sum => CSA_sum_2_29_2, c_out => CSA_carry_2_29_2);
FA_lbl_2_29_3: FA port map(in1 => CSA_carry_1_28_2, in2 => CSA_carry_1_28_1, c_in => CSA_carry_1_28_0, sum => CSA_sum_2_29_3, c_out => CSA_carry_2_29_3);
FA_lbl_2_30_0: FA port map(in1 => CSA_sum_1_30_6, in2 => CSA_sum_1_30_5, c_in => CSA_sum_1_30_4, sum => CSA_sum_2_30_0, c_out => CSA_carry_2_30_0);
FA_lbl_2_30_1: FA port map(in1 => CSA_sum_1_30_3, in2 => CSA_sum_1_30_2, c_in => CSA_sum_1_30_1, sum => CSA_sum_2_30_1, c_out => CSA_carry_2_30_1);
FA_lbl_2_30_2: FA port map(in1 => CSA_sum_1_30_0, in2 => CSA_carry_1_29_5, c_in => CSA_carry_1_29_4, sum => CSA_sum_2_30_2, c_out => CSA_carry_2_30_2);
FA_lbl_2_30_3: FA port map(in1 => CSA_carry_1_29_3, in2 => CSA_carry_1_29_2, c_in => CSA_carry_1_29_1, sum => CSA_sum_2_30_3, c_out => CSA_carry_2_30_3);
FA_lbl_2_31_0: FA port map(in1 => CSA_sum_1_31_6, in2 => CSA_sum_1_31_5, c_in => CSA_sum_1_31_4, sum => CSA_sum_2_31_0, c_out => CSA_carry_2_31_0);
FA_lbl_2_31_1: FA port map(in1 => CSA_sum_1_31_3, in2 => CSA_sum_1_31_2, c_in => CSA_sum_1_31_1, sum => CSA_sum_2_31_1, c_out => CSA_carry_2_31_1);
FA_lbl_2_31_2: FA port map(in1 => CSA_sum_1_31_0, in2 => CSA_carry_1_30_6, c_in => CSA_carry_1_30_5, sum => CSA_sum_2_31_2, c_out => CSA_carry_2_31_2);
FA_lbl_2_31_3: FA port map(in1 => CSA_carry_1_30_4, in2 => CSA_carry_1_30_3, c_in => CSA_carry_1_30_2, sum => CSA_sum_2_31_3, c_out => CSA_carry_2_31_3);
FA_lbl_2_31_4: FA port map(in1 => CSA_carry_1_30_1, in2 => CSA_carry_1_30_0, c_in => CSA_carry_0_30_0, sum => CSA_sum_2_31_4, c_out => CSA_carry_2_31_4);
FA_lbl_2_32_0: FA port map(in1 => CSA_sum_1_32_6, in2 => CSA_sum_1_32_5, c_in => CSA_sum_1_32_4, sum => CSA_sum_2_32_0, c_out => CSA_carry_2_32_0);
FA_lbl_2_32_1: FA port map(in1 => CSA_sum_1_32_3, in2 => CSA_sum_1_32_2, c_in => CSA_sum_1_32_1, sum => CSA_sum_2_32_1, c_out => CSA_carry_2_32_1);
FA_lbl_2_32_2: FA port map(in1 => CSA_sum_1_32_0, in2 => CSA_carry_1_31_6, c_in => CSA_carry_1_31_5, sum => CSA_sum_2_32_2, c_out => CSA_carry_2_32_2);
FA_lbl_2_32_3: FA port map(in1 => CSA_carry_1_31_4, in2 => CSA_carry_1_31_3, c_in => CSA_carry_1_31_2, sum => CSA_sum_2_32_3, c_out => CSA_carry_2_32_3);
FA_lbl_2_33_0: FA port map(in1 => CSA_sum_1_33_5, in2 => CSA_sum_1_33_4, c_in => CSA_sum_1_33_3, sum => CSA_sum_2_33_0, c_out => CSA_carry_2_33_0);
FA_lbl_2_33_1: FA port map(in1 => CSA_sum_1_33_2, in2 => CSA_sum_1_33_1, c_in => CSA_sum_1_33_0, sum => CSA_sum_2_33_1, c_out => CSA_carry_2_33_1);
FA_lbl_2_33_2: FA port map(in1 => CSA_carry_1_32_6, in2 => CSA_carry_1_32_5, c_in => CSA_carry_1_32_4, sum => CSA_sum_2_33_2, c_out => CSA_carry_2_33_2);
FA_lbl_2_33_3: FA port map(in1 => CSA_carry_1_32_3, in2 => CSA_carry_1_32_2, c_in => CSA_carry_1_32_1, sum => CSA_sum_2_33_3, c_out => CSA_carry_2_33_3);
FA_lbl_2_33_4: FA port map(in1 => CSA_carry_1_32_0, in2 => CSA_carry_0_32_1, c_in => CSA_carry_0_32_0, sum => CSA_sum_2_33_4, c_out => CSA_carry_2_33_4);
FA_lbl_2_34_0: FA port map(in1 => CSA_sum_1_34_6, in2 => CSA_sum_1_34_5, c_in => CSA_sum_1_34_4, sum => CSA_sum_2_34_0, c_out => CSA_carry_2_34_0);
FA_lbl_2_34_1: FA port map(in1 => CSA_sum_1_34_3, in2 => CSA_sum_1_34_2, c_in => CSA_sum_1_34_1, sum => CSA_sum_2_34_1, c_out => CSA_carry_2_34_1);
FA_lbl_2_34_2: FA port map(in1 => CSA_sum_1_34_0, in2 => CSA_carry_1_33_5, c_in => CSA_carry_1_33_4, sum => CSA_sum_2_34_2, c_out => CSA_carry_2_34_2);
FA_lbl_2_34_3: FA port map(in1 => CSA_carry_1_33_3, in2 => CSA_carry_1_33_2, c_in => CSA_carry_1_33_1, sum => CSA_sum_2_34_3, c_out => CSA_carry_2_34_3);
FA_lbl_2_35_0: FA port map(in1 => CSA_sum_1_35_5, in2 => CSA_sum_1_35_4, c_in => CSA_sum_1_35_3, sum => CSA_sum_2_35_0, c_out => CSA_carry_2_35_0);
FA_lbl_2_35_1: FA port map(in1 => CSA_sum_1_35_2, in2 => CSA_sum_1_35_1, c_in => CSA_sum_1_35_0, sum => CSA_sum_2_35_1, c_out => CSA_carry_2_35_1);
FA_lbl_2_35_2: FA port map(in1 => CSA_carry_1_34_6, in2 => CSA_carry_1_34_5, c_in => CSA_carry_1_34_4, sum => CSA_sum_2_35_2, c_out => CSA_carry_2_35_2);
FA_lbl_2_35_3: FA port map(in1 => CSA_carry_1_34_3, in2 => CSA_carry_1_34_2, c_in => CSA_carry_1_34_1, sum => CSA_sum_2_35_3, c_out => CSA_carry_2_35_3);
FA_lbl_2_36_0: FA port map(in1 => CSA_sum_1_36_5, in2 => CSA_sum_1_36_4, c_in => CSA_sum_1_36_3, sum => CSA_sum_2_36_0, c_out => CSA_carry_2_36_0);
FA_lbl_2_36_1: FA port map(in1 => CSA_sum_1_36_2, in2 => CSA_sum_1_36_1, c_in => CSA_sum_1_36_0, sum => CSA_sum_2_36_1, c_out => CSA_carry_2_36_1);
FA_lbl_2_36_2: FA port map(in1 => CSA_carry_1_35_5, in2 => CSA_carry_1_35_4, c_in => CSA_carry_1_35_3, sum => CSA_sum_2_36_2, c_out => CSA_carry_2_36_2);
FA_lbl_2_36_3: FA port map(in1 => CSA_carry_1_35_2, in2 => CSA_carry_1_35_1, c_in => CSA_carry_1_35_0, sum => CSA_sum_2_36_3, c_out => CSA_carry_2_36_3);
FA_lbl_2_37_0: FA port map(in1 => CSA_sum_1_37_5, in2 => CSA_sum_1_37_4, c_in => CSA_sum_1_37_3, sum => CSA_sum_2_37_0, c_out => CSA_carry_2_37_0);
FA_lbl_2_37_1: FA port map(in1 => CSA_sum_1_37_2, in2 => CSA_sum_1_37_1, c_in => CSA_sum_1_37_0, sum => CSA_sum_2_37_1, c_out => CSA_carry_2_37_1);
FA_lbl_2_37_2: FA port map(in1 => CSA_carry_1_36_5, in2 => CSA_carry_1_36_4, c_in => CSA_carry_1_36_3, sum => CSA_sum_2_37_2, c_out => CSA_carry_2_37_2);
FA_lbl_2_37_3: FA port map(in1 => CSA_carry_1_36_2, in2 => CSA_carry_1_36_1, c_in => CSA_carry_1_36_0, sum => CSA_sum_2_37_3, c_out => CSA_carry_2_37_3);
FA_lbl_2_38_0: FA port map(in1 => CSA_sum_1_38_4, in2 => CSA_sum_1_38_3, c_in => CSA_sum_1_38_2, sum => CSA_sum_2_38_0, c_out => CSA_carry_2_38_0);
FA_lbl_2_38_1: FA port map(in1 => CSA_sum_1_38_1, in2 => CSA_sum_1_38_0, c_in => CSA_carry_1_37_5, sum => CSA_sum_2_38_1, c_out => CSA_carry_2_38_1);
FA_lbl_2_38_2: FA port map(in1 => CSA_carry_1_37_4, in2 => CSA_carry_1_37_3, c_in => CSA_carry_1_37_2, sum => CSA_sum_2_38_2, c_out => CSA_carry_2_38_2);
FA_lbl_2_38_3: FA port map(in1 => CSA_carry_1_37_1, in2 => CSA_carry_1_37_0, c_in => CSA_carry_0_37_1, sum => CSA_sum_2_38_3, c_out => CSA_carry_2_38_3);
FA_lbl_2_39_0: FA port map(in1 => CSA_sum_1_39_4, in2 => CSA_sum_1_39_3, c_in => CSA_sum_1_39_2, sum => CSA_sum_2_39_0, c_out => CSA_carry_2_39_0);
FA_lbl_2_39_1: FA port map(in1 => CSA_sum_1_39_1, in2 => CSA_sum_1_39_0, c_in => CSA_carry_1_38_4, sum => CSA_sum_2_39_1, c_out => CSA_carry_2_39_1);
FA_lbl_2_39_2: FA port map(in1 => CSA_carry_1_38_3, in2 => CSA_carry_1_38_2, c_in => CSA_carry_1_38_1, sum => CSA_sum_2_39_2, c_out => CSA_carry_2_39_2);
FA_lbl_2_40_0: FA port map(in1 => CSA_sum_1_40_4, in2 => CSA_sum_1_40_3, c_in => CSA_sum_1_40_2, sum => CSA_sum_2_40_0, c_out => CSA_carry_2_40_0);
FA_lbl_2_40_1: FA port map(in1 => CSA_sum_1_40_1, in2 => CSA_sum_1_40_0, c_in => CSA_carry_1_39_4, sum => CSA_sum_2_40_1, c_out => CSA_carry_2_40_1);
FA_lbl_2_40_2: FA port map(in1 => CSA_carry_1_39_3, in2 => CSA_carry_1_39_2, c_in => CSA_carry_1_39_1, sum => CSA_sum_2_40_2, c_out => CSA_carry_2_40_2);
FA_lbl_2_40_3: FA port map(in1 => CSA_carry_1_39_0, in2 => CSA_carry_0_39_1, c_in => CSA_carry_0_39_0, sum => CSA_sum_2_40_3, c_out => CSA_carry_2_40_3);
FA_lbl_2_41_0: FA port map(in1 => CSA_sum_1_41_4, in2 => CSA_sum_1_41_3, c_in => CSA_sum_1_41_2, sum => CSA_sum_2_41_0, c_out => CSA_carry_2_41_0);
FA_lbl_2_41_1: FA port map(in1 => CSA_sum_1_41_1, in2 => CSA_sum_1_41_0, c_in => CSA_carry_1_40_4, sum => CSA_sum_2_41_1, c_out => CSA_carry_2_41_1);
FA_lbl_2_41_2: FA port map(in1 => CSA_carry_1_40_3, in2 => CSA_carry_1_40_2, c_in => CSA_carry_1_40_1, sum => CSA_sum_2_41_2, c_out => CSA_carry_2_41_2);
FA_lbl_2_42_0: FA port map(in1 => CSA_sum_1_42_3, in2 => CSA_sum_1_42_2, c_in => CSA_sum_1_42_1, sum => CSA_sum_2_42_0, c_out => CSA_carry_2_42_0);
FA_lbl_2_42_1: FA port map(in1 => CSA_sum_1_42_0, in2 => CSA_carry_1_41_4, c_in => CSA_carry_1_41_3, sum => CSA_sum_2_42_1, c_out => CSA_carry_2_42_1);
FA_lbl_2_42_2: FA port map(in1 => CSA_carry_1_41_2, in2 => CSA_carry_1_41_1, c_in => CSA_carry_1_41_0, sum => CSA_sum_2_42_2, c_out => CSA_carry_2_42_2);
FA_lbl_2_43_0: FA port map(in1 => CSA_sum_1_43_4, in2 => CSA_sum_1_43_3, c_in => CSA_sum_1_43_2, sum => CSA_sum_2_43_0, c_out => CSA_carry_2_43_0);
FA_lbl_2_43_1: FA port map(in1 => CSA_sum_1_43_1, in2 => CSA_sum_1_43_0, c_in => CSA_carry_1_42_3, sum => CSA_sum_2_43_1, c_out => CSA_carry_2_43_1);
FA_lbl_2_43_2: FA port map(in1 => CSA_carry_1_42_2, in2 => CSA_carry_1_42_1, c_in => CSA_carry_1_42_0, sum => CSA_sum_2_43_2, c_out => CSA_carry_2_43_2);
FA_lbl_2_44_0: FA port map(in1 => CSA_sum_1_44_3, in2 => CSA_sum_1_44_2, c_in => CSA_sum_1_44_1, sum => CSA_sum_2_44_0, c_out => CSA_carry_2_44_0);
FA_lbl_2_44_1: FA port map(in1 => CSA_sum_1_44_0, in2 => CSA_carry_1_43_4, c_in => CSA_carry_1_43_3, sum => CSA_sum_2_44_1, c_out => CSA_carry_2_44_1);
FA_lbl_2_44_2: FA port map(in1 => CSA_carry_1_43_2, in2 => CSA_carry_1_43_1, c_in => CSA_carry_1_43_0, sum => CSA_sum_2_44_2, c_out => CSA_carry_2_44_2);
FA_lbl_2_45_0: FA port map(in1 => CSA_sum_1_45_3, in2 => CSA_sum_1_45_2, c_in => CSA_sum_1_45_1, sum => CSA_sum_2_45_0, c_out => CSA_carry_2_45_0);
FA_lbl_2_45_1: FA port map(in1 => CSA_sum_1_45_0, in2 => CSA_carry_1_44_3, c_in => CSA_carry_1_44_2, sum => CSA_sum_2_45_1, c_out => CSA_carry_2_45_1);
FA_lbl_2_46_0: FA port map(in1 => CSA_sum_1_46_3, in2 => CSA_sum_1_46_2, c_in => CSA_sum_1_46_1, sum => CSA_sum_2_46_0, c_out => CSA_carry_2_46_0);
FA_lbl_2_46_1: FA port map(in1 => CSA_sum_1_46_0, in2 => CSA_carry_1_45_3, c_in => CSA_carry_1_45_2, sum => CSA_sum_2_46_1, c_out => CSA_carry_2_46_1);
FA_lbl_2_46_2: FA port map(in1 => CSA_carry_1_45_1, in2 => CSA_carry_1_45_0, c_in => CSA_carry_0_45_0, sum => CSA_sum_2_46_2, c_out => CSA_carry_2_46_2);
FA_lbl_2_47_0: FA port map(in1 => CSA_sum_1_47_2, in2 => CSA_sum_1_47_1, c_in => CSA_sum_1_47_0, sum => CSA_sum_2_47_0, c_out => CSA_carry_2_47_0);
FA_lbl_2_47_1: FA port map(in1 => CSA_carry_1_46_3, in2 => CSA_carry_1_46_2, c_in => CSA_carry_1_46_1, sum => CSA_sum_2_47_1, c_out => CSA_carry_2_47_1);
FA_lbl_2_47_2: FA port map(in1 => CSA_carry_1_46_0, in2 => CSA_carry_0_46_1, c_in => CSA_carry_0_46_0, sum => CSA_sum_2_47_2, c_out => CSA_carry_2_47_2);
FA_lbl_2_48_0: FA port map(in1 => CSA_sum_1_48_2, in2 => CSA_sum_1_48_1, c_in => CSA_sum_1_48_0, sum => CSA_sum_2_48_0, c_out => CSA_carry_2_48_0);
FA_lbl_2_48_1: FA port map(in1 => CSA_carry_1_47_2, in2 => CSA_carry_1_47_1, c_in => CSA_carry_1_47_0, sum => CSA_sum_2_48_1, c_out => CSA_carry_2_48_1);
FA_lbl_2_49_0: FA port map(in1 => CSA_sum_1_49_2, in2 => CSA_sum_1_49_1, c_in => CSA_sum_1_49_0, sum => CSA_sum_2_49_0, c_out => CSA_carry_2_49_0);
FA_lbl_2_49_1: FA port map(in1 => CSA_carry_1_48_2, in2 => CSA_carry_1_48_1, c_in => CSA_carry_1_48_0, sum => CSA_sum_2_49_1, c_out => CSA_carry_2_49_1);
FA_lbl_2_50_0: FA port map(in1 => CSA_sum_1_50_2, in2 => CSA_sum_1_50_1, c_in => CSA_sum_1_50_0, sum => CSA_sum_2_50_0, c_out => CSA_carry_2_50_0);
FA_lbl_2_50_1: FA port map(in1 => CSA_carry_1_49_2, in2 => CSA_carry_1_49_1, c_in => CSA_carry_1_49_0, sum => CSA_sum_2_50_1, c_out => CSA_carry_2_50_1);
FA_lbl_2_51_0: FA port map(in1 => CSA_sum_1_51_1, in2 => CSA_sum_1_51_0, c_in => CSA_carry_1_50_2, sum => CSA_sum_2_51_0, c_out => CSA_carry_2_51_0);
FA_lbl_2_51_1: FA port map(in1 => CSA_carry_1_50_1, in2 => CSA_carry_1_50_0, c_in => CSA_carry_0_50_1, sum => CSA_sum_2_51_1, c_out => CSA_carry_2_51_1);
FA_lbl_2_52_0: FA port map(in1 => CSA_sum_1_52_2, in2 => CSA_sum_1_52_1, c_in => CSA_sum_1_52_0, sum => CSA_sum_2_52_0, c_out => CSA_carry_2_52_0);
FA_lbl_2_53_0: FA port map(in1 => CSA_sum_1_53_1, in2 => CSA_sum_1_53_0, c_in => CSA_carry_1_52_2, sum => CSA_sum_2_53_0, c_out => CSA_carry_2_53_0);
FA_lbl_2_53_1: FA port map(in1 => CSA_carry_1_52_1, in2 => CSA_carry_1_52_0, c_in => CSA_carry_0_52_0, sum => CSA_sum_2_53_1, c_out => CSA_carry_2_53_1);
FA_lbl_2_54_0: FA port map(in1 => CSA_sum_1_54_1, in2 => CSA_sum_1_54_0, c_in => CSA_carry_1_53_1, sum => CSA_sum_2_54_0, c_out => CSA_carry_2_54_0);
FA_lbl_2_55_0: FA port map(in1 => CSA_sum_1_55_1, in2 => CSA_sum_1_55_0, c_in => CSA_carry_1_54_1, sum => CSA_sum_2_55_0, c_out => CSA_carry_2_55_0);
FA_lbl_2_56_0: FA port map(in1 => CSA_sum_1_56_0, in2 => CSA_carry_1_55_1, c_in => CSA_carry_1_55_0, sum => CSA_sum_2_56_0, c_out => CSA_carry_2_56_0);
FA_lbl_2_57_0: FA port map(in1 => CSA_sum_1_57_0, in2 => CSA_carry_1_56_0, c_in => CSA_carry_0_56_0, sum => CSA_sum_2_57_0, c_out => CSA_carry_2_57_0);
FA_lbl_2_58_0: FA port map(in1 => CSA_sum_1_58_0, in2 => CSA_carry_1_57_0, c_in => CSA_carry_0_57_1, sum => CSA_sum_2_58_0, c_out => CSA_carry_2_58_0);
FA_lbl_2_60_0: FA port map(in1 => CSA_carry_1_59_0, in2 => CSA_sum_0_60_0, c_in => CSA_carry_0_59_0, sum => CSA_sum_2_60_0, c_out => CSA_carry_2_60_0);
FA_lbl_3_5_0: FA port map(in1 => CSA_carry_2_4_0, in2 => CSA_sum_1_5_0, c_in => CSA_carry_1_4_0, sum => CSA_sum_3_5_0, c_out => CSA_carry_3_5_0);
FA_lbl_3_8_0: FA port map(in1 => CSA_sum_2_8_0, in2 => CSA_carry_2_7_0, c_in => CSA_carry_0_7_1, sum => CSA_sum_3_8_0, c_out => CSA_carry_3_8_0);
FA_lbl_3_9_0: FA port map(in1 => CSA_sum_2_9_0, in2 => CSA_carry_2_8_0, c_in => CSA_carry_0_8_0, sum => CSA_sum_3_9_0, c_out => CSA_carry_3_9_0);
FA_lbl_3_10_0: FA port map(in1 => CSA_sum_2_10_1, in2 => CSA_sum_2_10_0, c_in => CSA_carry_2_9_0, sum => CSA_sum_3_10_0, c_out => CSA_carry_3_10_0);
FA_lbl_3_11_0: FA port map(in1 => CSA_sum_2_11_0, in2 => CSA_carry_2_10_1, c_in => CSA_carry_2_10_0, sum => CSA_sum_3_11_0, c_out => CSA_carry_3_11_0);
FA_lbl_3_12_0: FA port map(in1 => CSA_sum_2_12_0, in2 => CSA_carry_2_11_0, c_in => CSA_carry_1_11_1, sum => CSA_sum_3_12_0, c_out => CSA_carry_3_12_0);
FA_lbl_3_13_0: FA port map(in1 => CSA_sum_2_13_1, in2 => CSA_sum_2_13_0, c_in => CSA_carry_2_12_0, sum => CSA_sum_3_13_0, c_out => CSA_carry_3_13_0);
FA_lbl_3_14_0: FA port map(in1 => CSA_sum_2_14_1, in2 => CSA_sum_2_14_0, c_in => CSA_carry_2_13_1, sum => CSA_sum_3_14_0, c_out => CSA_carry_3_14_0);
FA_lbl_3_15_0: FA port map(in1 => CSA_sum_2_15_1, in2 => CSA_sum_2_15_0, c_in => CSA_carry_2_14_1, sum => CSA_sum_3_15_0, c_out => CSA_carry_3_15_0);
FA_lbl_3_15_1: FA port map(in1 => CSA_carry_2_14_0, in2 => CSA_carry_0_14_1, c_in => CSA_carry_0_14_0, sum => CSA_sum_3_15_1, c_out => CSA_carry_3_15_1);
FA_lbl_3_16_0: FA port map(in1 => CSA_sum_2_16_1, in2 => CSA_sum_2_16_0, c_in => CSA_carry_2_15_1, sum => CSA_sum_3_16_0, c_out => CSA_carry_3_16_0);
FA_lbl_3_17_0: FA port map(in1 => CSA_sum_2_17_2, in2 => CSA_sum_2_17_1, c_in => CSA_sum_2_17_0, sum => CSA_sum_3_17_0, c_out => CSA_carry_3_17_0);
FA_lbl_3_18_0: FA port map(in1 => CSA_sum_2_18_1, in2 => CSA_sum_2_18_0, c_in => CSA_carry_2_17_2, sum => CSA_sum_3_18_0, c_out => CSA_carry_3_18_0);
FA_lbl_3_18_1: FA port map(in1 => CSA_carry_2_17_1, in2 => CSA_carry_2_17_0, c_in => CSA_carry_1_17_0, sum => CSA_sum_3_18_1, c_out => CSA_carry_3_18_1);
FA_lbl_3_19_0: FA port map(in1 => CSA_sum_2_19_2, in2 => CSA_sum_2_19_1, c_in => CSA_sum_2_19_0, sum => CSA_sum_3_19_0, c_out => CSA_carry_3_19_0);
FA_lbl_3_19_1: FA port map(in1 => CSA_carry_2_18_1, in2 => CSA_carry_2_18_0, c_in => CSA_carry_0_18_0, sum => CSA_sum_3_19_1, c_out => CSA_carry_3_19_1);
FA_lbl_3_20_0: FA port map(in1 => CSA_sum_2_20_2, in2 => CSA_sum_2_20_1, c_in => CSA_sum_2_20_0, sum => CSA_sum_3_20_0, c_out => CSA_carry_3_20_0);
FA_lbl_3_20_1: FA port map(in1 => CSA_carry_2_19_2, in2 => CSA_carry_2_19_1, c_in => CSA_carry_2_19_0, sum => CSA_sum_3_20_1, c_out => CSA_carry_3_20_1);
FA_lbl_3_21_0: FA port map(in1 => CSA_sum_2_21_2, in2 => CSA_sum_2_21_1, c_in => CSA_sum_2_21_0, sum => CSA_sum_3_21_0, c_out => CSA_carry_3_21_0);
FA_lbl_3_21_1: FA port map(in1 => CSA_carry_2_20_2, in2 => CSA_carry_2_20_1, c_in => CSA_carry_2_20_0, sum => CSA_sum_3_21_1, c_out => CSA_carry_3_21_1);
FA_lbl_3_22_0: FA port map(in1 => CSA_sum_2_22_2, in2 => CSA_sum_2_22_1, c_in => CSA_sum_2_22_0, sum => CSA_sum_3_22_0, c_out => CSA_carry_3_22_0);
FA_lbl_3_22_1: FA port map(in1 => CSA_carry_2_21_2, in2 => CSA_carry_2_21_1, c_in => CSA_carry_2_21_0, sum => CSA_sum_3_22_1, c_out => CSA_carry_3_22_1);
FA_lbl_3_23_0: FA port map(in1 => CSA_sum_2_23_2, in2 => CSA_sum_2_23_1, c_in => CSA_sum_2_23_0, sum => CSA_sum_3_23_0, c_out => CSA_carry_3_23_0);
FA_lbl_3_23_1: FA port map(in1 => CSA_carry_2_22_2, in2 => CSA_carry_2_22_1, c_in => CSA_carry_2_22_0, sum => CSA_sum_3_23_1, c_out => CSA_carry_3_23_1);
FA_lbl_3_24_0: FA port map(in1 => CSA_sum_2_24_3, in2 => CSA_sum_2_24_2, c_in => CSA_sum_2_24_1, sum => CSA_sum_3_24_0, c_out => CSA_carry_3_24_0);
FA_lbl_3_24_1: FA port map(in1 => CSA_sum_2_24_0, in2 => CSA_carry_2_23_2, c_in => CSA_carry_2_23_1, sum => CSA_sum_3_24_1, c_out => CSA_carry_3_24_1);
FA_lbl_3_25_0: FA port map(in1 => CSA_sum_2_25_2, in2 => CSA_sum_2_25_1, c_in => CSA_sum_2_25_0, sum => CSA_sum_3_25_0, c_out => CSA_carry_3_25_0);
FA_lbl_3_25_1: FA port map(in1 => CSA_carry_2_24_3, in2 => CSA_carry_2_24_2, c_in => CSA_carry_2_24_1, sum => CSA_sum_3_25_1, c_out => CSA_carry_3_25_1);
FA_lbl_3_25_2: FA port map(in1 => CSA_carry_2_24_0, in2 => CSA_carry_1_24_1, c_in => CSA_carry_1_24_0, sum => CSA_sum_3_25_2, c_out => CSA_carry_3_25_2);
FA_lbl_3_26_0: FA port map(in1 => CSA_sum_2_26_3, in2 => CSA_sum_2_26_2, c_in => CSA_sum_2_26_1, sum => CSA_sum_3_26_0, c_out => CSA_carry_3_26_0);
FA_lbl_3_26_1: FA port map(in1 => CSA_sum_2_26_0, in2 => CSA_carry_2_25_2, c_in => CSA_carry_2_25_1, sum => CSA_sum_3_26_1, c_out => CSA_carry_3_26_1);
FA_lbl_3_27_0: FA port map(in1 => CSA_sum_2_27_3, in2 => CSA_sum_2_27_2, c_in => CSA_sum_2_27_1, sum => CSA_sum_3_27_0, c_out => CSA_carry_3_27_0);
FA_lbl_3_27_1: FA port map(in1 => CSA_sum_2_27_0, in2 => CSA_carry_2_26_3, c_in => CSA_carry_2_26_2, sum => CSA_sum_3_27_1, c_out => CSA_carry_3_27_1);
FA_lbl_3_28_0: FA port map(in1 => CSA_sum_2_28_3, in2 => CSA_sum_2_28_2, c_in => CSA_sum_2_28_1, sum => CSA_sum_3_28_0, c_out => CSA_carry_3_28_0);
FA_lbl_3_28_1: FA port map(in1 => CSA_sum_2_28_0, in2 => CSA_carry_2_27_3, c_in => CSA_carry_2_27_2, sum => CSA_sum_3_28_1, c_out => CSA_carry_3_28_1);
FA_lbl_3_28_2: FA port map(in1 => CSA_carry_2_27_1, in2 => CSA_carry_2_27_0, c_in => CSA_carry_0_27_1, sum => CSA_sum_3_28_2, c_out => CSA_carry_3_28_2);
FA_lbl_3_29_0: FA port map(in1 => CSA_sum_2_29_3, in2 => CSA_sum_2_29_2, c_in => CSA_sum_2_29_1, sum => CSA_sum_3_29_0, c_out => CSA_carry_3_29_0);
FA_lbl_3_29_1: FA port map(in1 => CSA_sum_2_29_0, in2 => CSA_carry_2_28_3, c_in => CSA_carry_2_28_2, sum => CSA_sum_3_29_1, c_out => CSA_carry_3_29_1);
FA_lbl_3_29_2: FA port map(in1 => CSA_carry_2_28_1, in2 => CSA_carry_2_28_0, c_in => CSA_carry_0_28_0, sum => CSA_sum_3_29_2, c_out => CSA_carry_3_29_2);
FA_lbl_3_30_0: FA port map(in1 => CSA_sum_2_30_3, in2 => CSA_sum_2_30_2, c_in => CSA_sum_2_30_1, sum => CSA_sum_3_30_0, c_out => CSA_carry_3_30_0);
FA_lbl_3_30_1: FA port map(in1 => CSA_sum_2_30_0, in2 => CSA_carry_2_29_3, c_in => CSA_carry_2_29_2, sum => CSA_sum_3_30_1, c_out => CSA_carry_3_30_1);
FA_lbl_3_30_2: FA port map(in1 => CSA_carry_2_29_1, in2 => CSA_carry_2_29_0, c_in => CSA_carry_1_29_0, sum => CSA_sum_3_30_2, c_out => CSA_carry_3_30_2);
FA_lbl_3_31_0: FA port map(in1 => CSA_sum_2_31_4, in2 => CSA_sum_2_31_3, c_in => CSA_sum_2_31_2, sum => CSA_sum_3_31_0, c_out => CSA_carry_3_31_0);
FA_lbl_3_31_1: FA port map(in1 => CSA_sum_2_31_1, in2 => CSA_sum_2_31_0, c_in => CSA_carry_2_30_3, sum => CSA_sum_3_31_1, c_out => CSA_carry_3_31_1);
FA_lbl_3_31_2: FA port map(in1 => CSA_carry_2_30_2, in2 => CSA_carry_2_30_1, c_in => CSA_carry_2_30_0, sum => CSA_sum_3_31_2, c_out => CSA_carry_3_31_2);
FA_lbl_3_32_0: FA port map(in1 => CSA_sum_2_32_3, in2 => CSA_sum_2_32_2, c_in => CSA_sum_2_32_1, sum => CSA_sum_3_32_0, c_out => CSA_carry_3_32_0);
FA_lbl_3_32_1: FA port map(in1 => CSA_sum_2_32_0, in2 => CSA_carry_2_31_4, c_in => CSA_carry_2_31_3, sum => CSA_sum_3_32_1, c_out => CSA_carry_3_32_1);
FA_lbl_3_32_2: FA port map(in1 => CSA_carry_2_31_2, in2 => CSA_carry_2_31_1, c_in => CSA_carry_2_31_0, sum => CSA_sum_3_32_2, c_out => CSA_carry_3_32_2);
FA_lbl_3_33_0: FA port map(in1 => CSA_sum_2_33_4, in2 => CSA_sum_2_33_3, c_in => CSA_sum_2_33_2, sum => CSA_sum_3_33_0, c_out => CSA_carry_3_33_0);
FA_lbl_3_33_1: FA port map(in1 => CSA_sum_2_33_1, in2 => CSA_sum_2_33_0, c_in => CSA_carry_2_32_3, sum => CSA_sum_3_33_1, c_out => CSA_carry_3_33_1);
FA_lbl_3_33_2: FA port map(in1 => CSA_carry_2_32_2, in2 => CSA_carry_2_32_1, c_in => CSA_carry_2_32_0, sum => CSA_sum_3_33_2, c_out => CSA_carry_3_33_2);
FA_lbl_3_34_0: FA port map(in1 => CSA_sum_2_34_3, in2 => CSA_sum_2_34_2, c_in => CSA_sum_2_34_1, sum => CSA_sum_3_34_0, c_out => CSA_carry_3_34_0);
FA_lbl_3_34_1: FA port map(in1 => CSA_sum_2_34_0, in2 => CSA_carry_2_33_4, c_in => CSA_carry_2_33_3, sum => CSA_sum_3_34_1, c_out => CSA_carry_3_34_1);
FA_lbl_3_34_2: FA port map(in1 => CSA_carry_2_33_2, in2 => CSA_carry_2_33_1, c_in => CSA_carry_2_33_0, sum => CSA_sum_3_34_2, c_out => CSA_carry_3_34_2);
FA_lbl_3_35_0: FA port map(in1 => CSA_sum_2_35_3, in2 => CSA_sum_2_35_2, c_in => CSA_sum_2_35_1, sum => CSA_sum_3_35_0, c_out => CSA_carry_3_35_0);
FA_lbl_3_35_1: FA port map(in1 => CSA_sum_2_35_0, in2 => CSA_carry_2_34_3, c_in => CSA_carry_2_34_2, sum => CSA_sum_3_35_1, c_out => CSA_carry_3_35_1);
FA_lbl_3_35_2: FA port map(in1 => CSA_carry_2_34_1, in2 => CSA_carry_2_34_0, c_in => CSA_carry_1_34_0, sum => CSA_sum_3_35_2, c_out => CSA_carry_3_35_2);
FA_lbl_3_36_0: FA port map(in1 => CSA_sum_2_36_3, in2 => CSA_sum_2_36_2, c_in => CSA_sum_2_36_1, sum => CSA_sum_3_36_0, c_out => CSA_carry_3_36_0);
FA_lbl_3_36_1: FA port map(in1 => CSA_sum_2_36_0, in2 => CSA_carry_2_35_3, c_in => CSA_carry_2_35_2, sum => CSA_sum_3_36_1, c_out => CSA_carry_3_36_1);
FA_lbl_3_37_0: FA port map(in1 => CSA_sum_2_37_3, in2 => CSA_sum_2_37_2, c_in => CSA_sum_2_37_1, sum => CSA_sum_3_37_0, c_out => CSA_carry_3_37_0);
FA_lbl_3_37_1: FA port map(in1 => CSA_sum_2_37_0, in2 => CSA_carry_2_36_3, c_in => CSA_carry_2_36_2, sum => CSA_sum_3_37_1, c_out => CSA_carry_3_37_1);
FA_lbl_3_37_2: FA port map(in1 => CSA_carry_2_36_1, in2 => CSA_carry_2_36_0, c_in => CSA_carry_0_36_0, sum => CSA_sum_3_37_2, c_out => CSA_carry_3_37_2);
FA_lbl_3_38_0: FA port map(in1 => CSA_sum_2_38_3, in2 => CSA_sum_2_38_2, c_in => CSA_sum_2_38_1, sum => CSA_sum_3_38_0, c_out => CSA_carry_3_38_0);
FA_lbl_3_38_1: FA port map(in1 => CSA_sum_2_38_0, in2 => CSA_carry_2_37_3, c_in => CSA_carry_2_37_2, sum => CSA_sum_3_38_1, c_out => CSA_carry_3_38_1);
FA_lbl_3_38_2: FA port map(in1 => CSA_carry_2_37_1, in2 => CSA_carry_2_37_0, c_in => CSA_carry_0_37_0, sum => CSA_sum_3_38_2, c_out => CSA_carry_3_38_2);
FA_lbl_3_39_0: FA port map(in1 => CSA_sum_2_39_2, in2 => CSA_sum_2_39_1, c_in => CSA_sum_2_39_0, sum => CSA_sum_3_39_0, c_out => CSA_carry_3_39_0);
FA_lbl_3_39_1: FA port map(in1 => CSA_carry_2_38_3, in2 => CSA_carry_2_38_2, c_in => CSA_carry_2_38_1, sum => CSA_sum_3_39_1, c_out => CSA_carry_3_39_1);
FA_lbl_3_39_2: FA port map(in1 => CSA_carry_2_38_0, in2 => CSA_carry_1_38_0, c_in => CSA_carry_0_38_0, sum => CSA_sum_3_39_2, c_out => CSA_carry_3_39_2);
FA_lbl_3_40_0: FA port map(in1 => CSA_sum_2_40_3, in2 => CSA_sum_2_40_2, c_in => CSA_sum_2_40_1, sum => CSA_sum_3_40_0, c_out => CSA_carry_3_40_0);
FA_lbl_3_40_1: FA port map(in1 => CSA_sum_2_40_0, in2 => CSA_carry_2_39_2, c_in => CSA_carry_2_39_1, sum => CSA_sum_3_40_1, c_out => CSA_carry_3_40_1);
FA_lbl_3_41_0: FA port map(in1 => CSA_sum_2_41_2, in2 => CSA_sum_2_41_1, c_in => CSA_sum_2_41_0, sum => CSA_sum_3_41_0, c_out => CSA_carry_3_41_0);
FA_lbl_3_41_1: FA port map(in1 => CSA_carry_2_40_3, in2 => CSA_carry_2_40_2, c_in => CSA_carry_2_40_1, sum => CSA_sum_3_41_1, c_out => CSA_carry_3_41_1);
FA_lbl_3_42_0: FA port map(in1 => CSA_sum_2_42_2, in2 => CSA_sum_2_42_1, c_in => CSA_sum_2_42_0, sum => CSA_sum_3_42_0, c_out => CSA_carry_3_42_0);
FA_lbl_3_42_1: FA port map(in1 => CSA_carry_2_41_2, in2 => CSA_carry_2_41_1, c_in => CSA_carry_2_41_0, sum => CSA_sum_3_42_1, c_out => CSA_carry_3_42_1);
FA_lbl_3_43_0: FA port map(in1 => CSA_sum_2_43_2, in2 => CSA_sum_2_43_1, c_in => CSA_sum_2_43_0, sum => CSA_sum_3_43_0, c_out => CSA_carry_3_43_0);
FA_lbl_3_43_1: FA port map(in1 => CSA_carry_2_42_2, in2 => CSA_carry_2_42_1, c_in => CSA_carry_2_42_0, sum => CSA_sum_3_43_1, c_out => CSA_carry_3_43_1);
FA_lbl_3_44_0: FA port map(in1 => CSA_sum_2_44_2, in2 => CSA_sum_2_44_1, c_in => CSA_sum_2_44_0, sum => CSA_sum_3_44_0, c_out => CSA_carry_3_44_0);
FA_lbl_3_44_1: FA port map(in1 => CSA_carry_2_43_2, in2 => CSA_carry_2_43_1, c_in => CSA_carry_2_43_0, sum => CSA_sum_3_44_1, c_out => CSA_carry_3_44_1);
FA_lbl_3_45_0: FA port map(in1 => CSA_sum_2_45_1, in2 => CSA_sum_2_45_0, c_in => CSA_carry_2_44_2, sum => CSA_sum_3_45_0, c_out => CSA_carry_3_45_0);
FA_lbl_3_45_1: FA port map(in1 => CSA_carry_2_44_1, in2 => CSA_carry_2_44_0, c_in => CSA_carry_1_44_1, sum => CSA_sum_3_45_1, c_out => CSA_carry_3_45_1);
FA_lbl_3_46_0: FA port map(in1 => CSA_sum_2_46_2, in2 => CSA_sum_2_46_1, c_in => CSA_sum_2_46_0, sum => CSA_sum_3_46_0, c_out => CSA_carry_3_46_0);
FA_lbl_3_47_0: FA port map(in1 => CSA_sum_2_47_2, in2 => CSA_sum_2_47_1, c_in => CSA_sum_2_47_0, sum => CSA_sum_3_47_0, c_out => CSA_carry_3_47_0);
FA_lbl_3_47_1: FA port map(in1 => CSA_carry_2_46_2, in2 => CSA_carry_2_46_1, c_in => CSA_carry_2_46_0, sum => CSA_sum_3_47_1, c_out => CSA_carry_3_47_1);
FA_lbl_3_48_0: FA port map(in1 => CSA_sum_2_48_1, in2 => CSA_sum_2_48_0, c_in => CSA_carry_2_47_2, sum => CSA_sum_3_48_0, c_out => CSA_carry_3_48_0);
FA_lbl_3_48_1: FA port map(in1 => CSA_carry_2_47_1, in2 => CSA_carry_2_47_0, c_in => CSA_carry_0_47_0, sum => CSA_sum_3_48_1, c_out => CSA_carry_3_48_1);
FA_lbl_3_49_0: FA port map(in1 => CSA_sum_2_49_1, in2 => CSA_sum_2_49_0, c_in => CSA_carry_2_48_1, sum => CSA_sum_3_49_0, c_out => CSA_carry_3_49_0);
FA_lbl_3_49_1: FA port map(in1 => CSA_carry_2_48_0, in2 => CSA_carry_0_48_1, c_in => CSA_carry_0_48_0, sum => CSA_sum_3_49_1, c_out => CSA_carry_3_49_1);
FA_lbl_3_50_0: FA port map(in1 => CSA_sum_2_50_1, in2 => CSA_sum_2_50_0, c_in => CSA_carry_2_49_1, sum => CSA_sum_3_50_0, c_out => CSA_carry_3_50_0);
FA_lbl_3_51_0: FA port map(in1 => CSA_sum_2_51_1, in2 => CSA_sum_2_51_0, c_in => CSA_carry_2_50_1, sum => CSA_sum_3_51_0, c_out => CSA_carry_3_51_0);
FA_lbl_3_52_0: FA port map(in1 => CSA_sum_2_52_0, in2 => CSA_carry_2_51_1, c_in => CSA_carry_2_51_0, sum => CSA_sum_3_52_0, c_out => CSA_carry_3_52_0);
FA_lbl_3_53_0: FA port map(in1 => CSA_sum_2_53_1, in2 => CSA_sum_2_53_0, c_in => CSA_carry_2_52_0, sum => CSA_sum_3_53_0, c_out => CSA_carry_3_53_0);
FA_lbl_3_54_0: FA port map(in1 => CSA_sum_2_54_0, in2 => CSA_carry_2_53_1, c_in => CSA_carry_2_53_0, sum => CSA_sum_3_54_0, c_out => CSA_carry_3_54_0);
FA_lbl_3_55_0: FA port map(in1 => CSA_sum_2_55_0, in2 => CSA_carry_2_54_0, c_in => CSA_carry_1_54_0, sum => CSA_sum_3_55_0, c_out => CSA_carry_3_55_0);
FA_lbl_3_56_0: FA port map(in1 => CSA_sum_2_56_0, in2 => CSA_carry_2_55_0, c_in => CSA_carry_0_55_1, sum => CSA_sum_3_56_0, c_out => CSA_carry_3_56_0);
FA_lbl_3_58_0: FA port map(in1 => CSA_sum_2_58_0, in2 => CSA_carry_2_57_0, c_in => CSA_carry_0_57_0, sum => CSA_sum_3_58_0, c_out => CSA_carry_3_58_0);
FA_lbl_3_59_0: FA port map(in1 => CSA_carry_2_58_0, in2 => CSA_sum_1_59_0, c_in => CSA_carry_1_58_0, sum => CSA_sum_3_59_0, c_out => CSA_carry_3_59_0);
FA_lbl_4_6_0: FA port map(in1 => CSA_carry_3_5_0, in2 => CSA_sum_2_6_0, c_in => CSA_carry_0_5_0, sum => CSA_sum_4_6_0, c_out => CSA_carry_4_6_0);
FA_lbl_4_11_0: FA port map(in1 => CSA_sum_3_11_0, in2 => CSA_carry_3_10_0, c_in => CSA_carry_1_10_0, sum => CSA_sum_4_11_0, c_out => CSA_carry_4_11_0);
FA_lbl_4_12_0: FA port map(in1 => CSA_sum_3_12_0, in2 => CSA_carry_3_11_0, c_in => CSA_carry_1_11_0, sum => CSA_sum_4_12_0, c_out => CSA_carry_4_12_0);
FA_lbl_4_13_0: FA port map(in1 => CSA_sum_3_13_0, in2 => CSA_carry_3_12_0, c_in => CSA_carry_0_12_0, sum => CSA_sum_4_13_0, c_out => CSA_carry_4_13_0);
FA_lbl_4_14_0: FA port map(in1 => CSA_sum_3_14_0, in2 => CSA_carry_3_13_0, c_in => CSA_carry_2_13_0, sum => CSA_sum_4_14_0, c_out => CSA_carry_4_14_0);
FA_lbl_4_15_0: FA port map(in1 => CSA_sum_3_15_1, in2 => CSA_sum_3_15_0, c_in => CSA_carry_3_14_0, sum => CSA_sum_4_15_0, c_out => CSA_carry_4_15_0);
FA_lbl_4_16_0: FA port map(in1 => CSA_sum_3_16_0, in2 => CSA_carry_3_15_1, c_in => CSA_carry_3_15_0, sum => CSA_sum_4_16_0, c_out => CSA_carry_4_16_0);
FA_lbl_4_17_0: FA port map(in1 => CSA_sum_3_17_0, in2 => CSA_carry_3_16_0, c_in => CSA_carry_2_16_1, sum => CSA_sum_4_17_0, c_out => CSA_carry_4_17_0);
FA_lbl_4_18_0: FA port map(in1 => CSA_sum_3_18_1, in2 => CSA_sum_3_18_0, c_in => CSA_carry_3_17_0, sum => CSA_sum_4_18_0, c_out => CSA_carry_4_18_0);
FA_lbl_4_19_0: FA port map(in1 => CSA_sum_3_19_1, in2 => CSA_sum_3_19_0, c_in => CSA_carry_3_18_1, sum => CSA_sum_4_19_0, c_out => CSA_carry_4_19_0);
FA_lbl_4_20_0: FA port map(in1 => CSA_sum_3_20_1, in2 => CSA_sum_3_20_0, c_in => CSA_carry_3_19_1, sum => CSA_sum_4_20_0, c_out => CSA_carry_4_20_0);
FA_lbl_4_21_0: FA port map(in1 => CSA_sum_3_21_1, in2 => CSA_sum_3_21_0, c_in => CSA_carry_3_20_1, sum => CSA_sum_4_21_0, c_out => CSA_carry_4_21_0);
FA_lbl_4_22_0: FA port map(in1 => CSA_sum_3_22_1, in2 => CSA_sum_3_22_0, c_in => CSA_carry_3_21_1, sum => CSA_sum_4_22_0, c_out => CSA_carry_4_22_0);
FA_lbl_4_22_1: FA port map(in1 => CSA_carry_3_21_0, in2 => CSA_carry_1_21_0, c_in => CSA_carry_0_21_0, sum => CSA_sum_4_22_1, c_out => CSA_carry_4_22_1);
FA_lbl_4_23_0: FA port map(in1 => CSA_sum_3_23_1, in2 => CSA_sum_3_23_0, c_in => CSA_carry_3_22_1, sum => CSA_sum_4_23_0, c_out => CSA_carry_4_23_0);
FA_lbl_4_24_0: FA port map(in1 => CSA_sum_3_24_1, in2 => CSA_sum_3_24_0, c_in => CSA_carry_3_23_1, sum => CSA_sum_4_24_0, c_out => CSA_carry_4_24_0);
FA_lbl_4_25_0: FA port map(in1 => CSA_sum_3_25_2, in2 => CSA_sum_3_25_1, c_in => CSA_sum_3_25_0, sum => CSA_sum_4_25_0, c_out => CSA_carry_4_25_0);
FA_lbl_4_26_0: FA port map(in1 => CSA_sum_3_26_1, in2 => CSA_sum_3_26_0, c_in => CSA_carry_3_25_2, sum => CSA_sum_4_26_0, c_out => CSA_carry_4_26_0);
FA_lbl_4_26_1: FA port map(in1 => CSA_carry_3_25_1, in2 => CSA_carry_3_25_0, c_in => CSA_carry_2_25_0, sum => CSA_sum_4_26_1, c_out => CSA_carry_4_26_1);
FA_lbl_4_27_0: FA port map(in1 => CSA_sum_3_27_1, in2 => CSA_sum_3_27_0, c_in => CSA_carry_3_26_1, sum => CSA_sum_4_27_0, c_out => CSA_carry_4_27_0);
FA_lbl_4_27_1: FA port map(in1 => CSA_carry_3_26_0, in2 => CSA_carry_2_26_1, c_in => CSA_carry_2_26_0, sum => CSA_sum_4_27_1, c_out => CSA_carry_4_27_1);
FA_lbl_4_28_0: FA port map(in1 => CSA_sum_3_28_2, in2 => CSA_sum_3_28_1, c_in => CSA_sum_3_28_0, sum => CSA_sum_4_28_0, c_out => CSA_carry_4_28_0);
FA_lbl_4_28_1: FA port map(in1 => CSA_carry_3_27_1, in2 => CSA_carry_3_27_0, c_in => CSA_carry_0_27_0, sum => CSA_sum_4_28_1, c_out => CSA_carry_4_28_1);
FA_lbl_4_29_0: FA port map(in1 => CSA_sum_3_29_2, in2 => CSA_sum_3_29_1, c_in => CSA_sum_3_29_0, sum => CSA_sum_4_29_0, c_out => CSA_carry_4_29_0);
FA_lbl_4_29_1: FA port map(in1 => CSA_carry_3_28_2, in2 => CSA_carry_3_28_1, c_in => CSA_carry_3_28_0, sum => CSA_sum_4_29_1, c_out => CSA_carry_4_29_1);
FA_lbl_4_30_0: FA port map(in1 => CSA_sum_3_30_2, in2 => CSA_sum_3_30_1, c_in => CSA_sum_3_30_0, sum => CSA_sum_4_30_0, c_out => CSA_carry_4_30_0);
FA_lbl_4_30_1: FA port map(in1 => CSA_carry_3_29_2, in2 => CSA_carry_3_29_1, c_in => CSA_carry_3_29_0, sum => CSA_sum_4_30_1, c_out => CSA_carry_4_30_1);
FA_lbl_4_31_0: FA port map(in1 => CSA_sum_3_31_2, in2 => CSA_sum_3_31_1, c_in => CSA_sum_3_31_0, sum => CSA_sum_4_31_0, c_out => CSA_carry_4_31_0);
FA_lbl_4_31_1: FA port map(in1 => CSA_carry_3_30_2, in2 => CSA_carry_3_30_1, c_in => CSA_carry_3_30_0, sum => CSA_sum_4_31_1, c_out => CSA_carry_4_31_1);
FA_lbl_4_32_0: FA port map(in1 => CSA_sum_3_32_2, in2 => CSA_sum_3_32_1, c_in => CSA_sum_3_32_0, sum => CSA_sum_4_32_0, c_out => CSA_carry_4_32_0);
FA_lbl_4_32_1: FA port map(in1 => CSA_carry_3_31_2, in2 => CSA_carry_3_31_1, c_in => CSA_carry_3_31_0, sum => CSA_sum_4_32_1, c_out => CSA_carry_4_32_1);
FA_lbl_4_33_0: FA port map(in1 => CSA_sum_3_33_2, in2 => CSA_sum_3_33_1, c_in => CSA_sum_3_33_0, sum => CSA_sum_4_33_0, c_out => CSA_carry_4_33_0);
FA_lbl_4_33_1: FA port map(in1 => CSA_carry_3_32_2, in2 => CSA_carry_3_32_1, c_in => CSA_carry_3_32_0, sum => CSA_sum_4_33_1, c_out => CSA_carry_4_33_1);
FA_lbl_4_34_0: FA port map(in1 => CSA_sum_3_34_2, in2 => CSA_sum_3_34_1, c_in => CSA_sum_3_34_0, sum => CSA_sum_4_34_0, c_out => CSA_carry_4_34_0);
FA_lbl_4_34_1: FA port map(in1 => CSA_carry_3_33_2, in2 => CSA_carry_3_33_1, c_in => CSA_carry_3_33_0, sum => CSA_sum_4_34_1, c_out => CSA_carry_4_34_1);
FA_lbl_4_35_0: FA port map(in1 => CSA_sum_3_35_2, in2 => CSA_sum_3_35_1, c_in => CSA_sum_3_35_0, sum => CSA_sum_4_35_0, c_out => CSA_carry_4_35_0);
FA_lbl_4_35_1: FA port map(in1 => CSA_carry_3_34_2, in2 => CSA_carry_3_34_1, c_in => CSA_carry_3_34_0, sum => CSA_sum_4_35_1, c_out => CSA_carry_4_35_1);
FA_lbl_4_36_0: FA port map(in1 => CSA_sum_3_36_1, in2 => CSA_sum_3_36_0, c_in => CSA_carry_3_35_2, sum => CSA_sum_4_36_0, c_out => CSA_carry_4_36_0);
FA_lbl_4_36_1: FA port map(in1 => CSA_carry_3_35_1, in2 => CSA_carry_3_35_0, c_in => CSA_carry_2_35_1, sum => CSA_sum_4_36_1, c_out => CSA_carry_4_36_1);
FA_lbl_4_37_0: FA port map(in1 => CSA_sum_3_37_2, in2 => CSA_sum_3_37_1, c_in => CSA_sum_3_37_0, sum => CSA_sum_4_37_0, c_out => CSA_carry_4_37_0);
FA_lbl_4_38_0: FA port map(in1 => CSA_sum_3_38_2, in2 => CSA_sum_3_38_1, c_in => CSA_sum_3_38_0, sum => CSA_sum_4_38_0, c_out => CSA_carry_4_38_0);
FA_lbl_4_38_1: FA port map(in1 => CSA_carry_3_37_2, in2 => CSA_carry_3_37_1, c_in => CSA_carry_3_37_0, sum => CSA_sum_4_38_1, c_out => CSA_carry_4_38_1);
FA_lbl_4_39_0: FA port map(in1 => CSA_sum_3_39_2, in2 => CSA_sum_3_39_1, c_in => CSA_sum_3_39_0, sum => CSA_sum_4_39_0, c_out => CSA_carry_4_39_0);
FA_lbl_4_39_1: FA port map(in1 => CSA_carry_3_38_2, in2 => CSA_carry_3_38_1, c_in => CSA_carry_3_38_0, sum => CSA_sum_4_39_1, c_out => CSA_carry_4_39_1);
FA_lbl_4_40_0: FA port map(in1 => CSA_sum_3_40_1, in2 => CSA_sum_3_40_0, c_in => CSA_carry_3_39_2, sum => CSA_sum_4_40_0, c_out => CSA_carry_4_40_0);
FA_lbl_4_40_1: FA port map(in1 => CSA_carry_3_39_1, in2 => CSA_carry_3_39_0, c_in => CSA_carry_2_39_0, sum => CSA_sum_4_40_1, c_out => CSA_carry_4_40_1);
FA_lbl_4_41_0: FA port map(in1 => CSA_sum_3_41_1, in2 => CSA_sum_3_41_0, c_in => CSA_carry_3_40_1, sum => CSA_sum_4_41_0, c_out => CSA_carry_4_41_0);
FA_lbl_4_41_1: FA port map(in1 => CSA_carry_3_40_0, in2 => CSA_carry_2_40_0, c_in => CSA_carry_1_40_0, sum => CSA_sum_4_41_1, c_out => CSA_carry_4_41_1);
FA_lbl_4_42_0: FA port map(in1 => CSA_sum_3_42_1, in2 => CSA_sum_3_42_0, c_in => CSA_carry_3_41_1, sum => CSA_sum_4_42_0, c_out => CSA_carry_4_42_0);
FA_lbl_4_42_1: FA port map(in1 => CSA_carry_3_41_0, in2 => CSA_carry_0_41_1, c_in => CSA_carry_0_41_0, sum => CSA_sum_4_42_1, c_out => CSA_carry_4_42_1);
FA_lbl_4_43_0: FA port map(in1 => CSA_sum_3_43_1, in2 => CSA_sum_3_43_0, c_in => CSA_carry_3_42_1, sum => CSA_sum_4_43_0, c_out => CSA_carry_4_43_0);
FA_lbl_4_44_0: FA port map(in1 => CSA_sum_3_44_1, in2 => CSA_sum_3_44_0, c_in => CSA_carry_3_43_1, sum => CSA_sum_4_44_0, c_out => CSA_carry_4_44_0);
FA_lbl_4_45_0: FA port map(in1 => CSA_sum_3_45_1, in2 => CSA_sum_3_45_0, c_in => CSA_carry_3_44_1, sum => CSA_sum_4_45_0, c_out => CSA_carry_4_45_0);
FA_lbl_4_46_0: FA port map(in1 => CSA_sum_3_46_0, in2 => CSA_carry_3_45_1, c_in => CSA_carry_3_45_0, sum => CSA_sum_4_46_0, c_out => CSA_carry_4_46_0);
FA_lbl_4_47_0: FA port map(in1 => CSA_sum_3_47_1, in2 => CSA_sum_3_47_0, c_in => CSA_carry_3_46_0, sum => CSA_sum_4_47_0, c_out => CSA_carry_4_47_0);
FA_lbl_4_48_0: FA port map(in1 => CSA_sum_3_48_1, in2 => CSA_sum_3_48_0, c_in => CSA_carry_3_47_1, sum => CSA_sum_4_48_0, c_out => CSA_carry_4_48_0);
FA_lbl_4_49_0: FA port map(in1 => CSA_sum_3_49_1, in2 => CSA_sum_3_49_0, c_in => CSA_carry_3_48_1, sum => CSA_sum_4_49_0, c_out => CSA_carry_4_49_0);
FA_lbl_4_50_0: FA port map(in1 => CSA_sum_3_50_0, in2 => CSA_carry_3_49_1, c_in => CSA_carry_3_49_0, sum => CSA_sum_4_50_0, c_out => CSA_carry_4_50_0);
FA_lbl_4_51_0: FA port map(in1 => CSA_sum_3_51_0, in2 => CSA_carry_3_50_0, c_in => CSA_carry_2_50_0, sum => CSA_sum_4_51_0, c_out => CSA_carry_4_51_0);
FA_lbl_4_52_0: FA port map(in1 => CSA_sum_3_52_0, in2 => CSA_carry_3_51_0, c_in => CSA_carry_1_51_1, sum => CSA_sum_4_52_0, c_out => CSA_carry_4_52_0);
FA_lbl_4_54_0: FA port map(in1 => CSA_sum_3_54_0, in2 => CSA_carry_3_53_0, c_in => CSA_carry_1_53_0, sum => CSA_sum_4_54_0, c_out => CSA_carry_4_54_0);
FA_lbl_4_55_0: FA port map(in1 => CSA_sum_3_55_0, in2 => CSA_carry_3_54_0, c_in => CSA_carry_0_54_0, sum => CSA_sum_4_55_0, c_out => CSA_carry_4_55_0);
FA_lbl_4_56_0: FA port map(in1 => CSA_sum_3_56_0, in2 => CSA_carry_3_55_0, c_in => CSA_carry_0_55_0, sum => CSA_sum_4_56_0, c_out => CSA_carry_4_56_0);
FA_lbl_4_57_0: FA port map(in1 => CSA_carry_3_56_0, in2 => CSA_sum_2_57_0, c_in => CSA_carry_2_56_0, sum => CSA_sum_4_57_0, c_out => CSA_carry_4_57_0);
FA_lbl_5_7_0: FA port map(in1 => CSA_carry_4_6_0, in2 => CSA_sum_2_7_0, c_in => CSA_carry_2_6_0, sum => CSA_sum_5_7_0, c_out => CSA_carry_5_7_0);
FA_lbl_5_16_0: FA port map(in1 => CSA_sum_4_16_0, in2 => CSA_carry_4_15_0, c_in => CSA_carry_2_15_0, sum => CSA_sum_5_16_0, c_out => CSA_carry_5_16_0);
FA_lbl_5_17_0: FA port map(in1 => CSA_sum_4_17_0, in2 => CSA_carry_4_16_0, c_in => CSA_carry_2_16_0, sum => CSA_sum_5_17_0, c_out => CSA_carry_5_17_0);
FA_lbl_5_18_0: FA port map(in1 => CSA_sum_4_18_0, in2 => CSA_carry_4_17_0, c_in => CSA_carry_0_17_0, sum => CSA_sum_5_18_0, c_out => CSA_carry_5_18_0);
FA_lbl_5_19_0: FA port map(in1 => CSA_sum_4_19_0, in2 => CSA_carry_4_18_0, c_in => CSA_carry_3_18_0, sum => CSA_sum_5_19_0, c_out => CSA_carry_5_19_0);
FA_lbl_5_20_0: FA port map(in1 => CSA_sum_4_20_0, in2 => CSA_carry_4_19_0, c_in => CSA_carry_3_19_0, sum => CSA_sum_5_20_0, c_out => CSA_carry_5_20_0);
FA_lbl_5_21_0: FA port map(in1 => CSA_sum_4_21_0, in2 => CSA_carry_4_20_0, c_in => CSA_carry_3_20_0, sum => CSA_sum_5_21_0, c_out => CSA_carry_5_21_0);
FA_lbl_5_22_0: FA port map(in1 => CSA_sum_4_22_1, in2 => CSA_sum_4_22_0, c_in => CSA_carry_4_21_0, sum => CSA_sum_5_22_0, c_out => CSA_carry_5_22_0);
FA_lbl_5_23_0: FA port map(in1 => CSA_sum_4_23_0, in2 => CSA_carry_4_22_1, c_in => CSA_carry_4_22_0, sum => CSA_sum_5_23_0, c_out => CSA_carry_5_23_0);
FA_lbl_5_24_0: FA port map(in1 => CSA_sum_4_24_0, in2 => CSA_carry_4_23_0, c_in => CSA_carry_3_23_0, sum => CSA_sum_5_24_0, c_out => CSA_carry_5_24_0);
FA_lbl_5_25_0: FA port map(in1 => CSA_sum_4_25_0, in2 => CSA_carry_4_24_0, c_in => CSA_carry_3_24_1, sum => CSA_sum_5_25_0, c_out => CSA_carry_5_25_0);
FA_lbl_5_26_0: FA port map(in1 => CSA_sum_4_26_1, in2 => CSA_sum_4_26_0, c_in => CSA_carry_4_25_0, sum => CSA_sum_5_26_0, c_out => CSA_carry_5_26_0);
FA_lbl_5_27_0: FA port map(in1 => CSA_sum_4_27_1, in2 => CSA_sum_4_27_0, c_in => CSA_carry_4_26_1, sum => CSA_sum_5_27_0, c_out => CSA_carry_5_27_0);
FA_lbl_5_28_0: FA port map(in1 => CSA_sum_4_28_1, in2 => CSA_sum_4_28_0, c_in => CSA_carry_4_27_1, sum => CSA_sum_5_28_0, c_out => CSA_carry_5_28_0);
FA_lbl_5_29_0: FA port map(in1 => CSA_sum_4_29_1, in2 => CSA_sum_4_29_0, c_in => CSA_carry_4_28_1, sum => CSA_sum_5_29_0, c_out => CSA_carry_5_29_0);
FA_lbl_5_30_0: FA port map(in1 => CSA_sum_4_30_1, in2 => CSA_sum_4_30_0, c_in => CSA_carry_4_29_1, sum => CSA_sum_5_30_0, c_out => CSA_carry_5_30_0);
FA_lbl_5_31_0: FA port map(in1 => CSA_sum_4_31_1, in2 => CSA_sum_4_31_0, c_in => CSA_carry_4_30_1, sum => CSA_sum_5_31_0, c_out => CSA_carry_5_31_0);
FA_lbl_5_32_0: FA port map(in1 => CSA_sum_4_32_1, in2 => CSA_sum_4_32_0, c_in => CSA_carry_4_31_1, sum => CSA_sum_5_32_0, c_out => CSA_carry_5_32_0);
FA_lbl_5_32_1: FA port map(in1 => CSA_carry_4_31_0, in2 => CSA_carry_1_31_1, c_in => CSA_carry_1_31_0, sum => CSA_sum_5_32_1, c_out => CSA_carry_5_32_1);
FA_lbl_5_33_0: FA port map(in1 => CSA_sum_4_33_1, in2 => CSA_sum_4_33_0, c_in => CSA_carry_4_32_1, sum => CSA_sum_5_33_0, c_out => CSA_carry_5_33_0);
FA_lbl_5_34_0: FA port map(in1 => CSA_sum_4_34_1, in2 => CSA_sum_4_34_0, c_in => CSA_carry_4_33_1, sum => CSA_sum_5_34_0, c_out => CSA_carry_5_34_0);
FA_lbl_5_35_0: FA port map(in1 => CSA_sum_4_35_1, in2 => CSA_sum_4_35_0, c_in => CSA_carry_4_34_1, sum => CSA_sum_5_35_0, c_out => CSA_carry_5_35_0);
FA_lbl_5_36_0: FA port map(in1 => CSA_sum_4_36_1, in2 => CSA_sum_4_36_0, c_in => CSA_carry_4_35_1, sum => CSA_sum_5_36_0, c_out => CSA_carry_5_36_0);
FA_lbl_5_37_0: FA port map(in1 => CSA_sum_4_37_0, in2 => CSA_carry_4_36_1, c_in => CSA_carry_4_36_0, sum => CSA_sum_5_37_0, c_out => CSA_carry_5_37_0);
FA_lbl_5_38_0: FA port map(in1 => CSA_sum_4_38_1, in2 => CSA_sum_4_38_0, c_in => CSA_carry_4_37_0, sum => CSA_sum_5_38_0, c_out => CSA_carry_5_38_0);
FA_lbl_5_39_0: FA port map(in1 => CSA_sum_4_39_1, in2 => CSA_sum_4_39_0, c_in => CSA_carry_4_38_1, sum => CSA_sum_5_39_0, c_out => CSA_carry_5_39_0);
FA_lbl_5_40_0: FA port map(in1 => CSA_sum_4_40_1, in2 => CSA_sum_4_40_0, c_in => CSA_carry_4_39_1, sum => CSA_sum_5_40_0, c_out => CSA_carry_5_40_0);
FA_lbl_5_41_0: FA port map(in1 => CSA_sum_4_41_1, in2 => CSA_sum_4_41_0, c_in => CSA_carry_4_40_1, sum => CSA_sum_5_41_0, c_out => CSA_carry_5_41_0);
FA_lbl_5_42_0: FA port map(in1 => CSA_sum_4_42_1, in2 => CSA_sum_4_42_0, c_in => CSA_carry_4_41_1, sum => CSA_sum_5_42_0, c_out => CSA_carry_5_42_0);
FA_lbl_5_43_0: FA port map(in1 => CSA_sum_4_43_0, in2 => CSA_carry_4_42_1, c_in => CSA_carry_4_42_0, sum => CSA_sum_5_43_0, c_out => CSA_carry_5_43_0);
FA_lbl_5_44_0: FA port map(in1 => CSA_sum_4_44_0, in2 => CSA_carry_4_43_0, c_in => CSA_carry_3_43_0, sum => CSA_sum_5_44_0, c_out => CSA_carry_5_44_0);
FA_lbl_5_45_0: FA port map(in1 => CSA_sum_4_45_0, in2 => CSA_carry_4_44_0, c_in => CSA_carry_3_44_0, sum => CSA_sum_5_45_0, c_out => CSA_carry_5_45_0);
FA_lbl_5_46_0: FA port map(in1 => CSA_sum_4_46_0, in2 => CSA_carry_4_45_0, c_in => CSA_carry_2_45_1, sum => CSA_sum_5_46_0, c_out => CSA_carry_5_46_0);
FA_lbl_5_48_0: FA port map(in1 => CSA_sum_4_48_0, in2 => CSA_carry_4_47_0, c_in => CSA_carry_3_47_0, sum => CSA_sum_5_48_0, c_out => CSA_carry_5_48_0);
FA_lbl_5_49_0: FA port map(in1 => CSA_sum_4_49_0, in2 => CSA_carry_4_48_0, c_in => CSA_carry_3_48_0, sum => CSA_sum_5_49_0, c_out => CSA_carry_5_49_0);
FA_lbl_5_50_0: FA port map(in1 => CSA_sum_4_50_0, in2 => CSA_carry_4_49_0, c_in => CSA_carry_2_49_0, sum => CSA_sum_5_50_0, c_out => CSA_carry_5_50_0);
FA_lbl_5_51_0: FA port map(in1 => CSA_sum_4_51_0, in2 => CSA_carry_4_50_0, c_in => CSA_carry_0_50_0, sum => CSA_sum_5_51_0, c_out => CSA_carry_5_51_0);
FA_lbl_5_52_0: FA port map(in1 => CSA_sum_4_52_0, in2 => CSA_carry_4_51_0, c_in => CSA_carry_1_51_0, sum => CSA_sum_5_52_0, c_out => CSA_carry_5_52_0);
FA_lbl_5_53_0: FA port map(in1 => CSA_carry_4_52_0, in2 => CSA_sum_3_53_0, c_in => CSA_carry_3_52_0, sum => CSA_sum_5_53_0, c_out => CSA_carry_5_53_0);
FA_lbl_6_8_0: FA port map(in1 => CSA_carry_5_7_0, in2 => CSA_sum_3_8_0, c_in => CSA_carry_0_7_0, sum => CSA_sum_6_8_0, c_out => CSA_carry_6_8_0);
FA_lbl_6_23_0: FA port map(in1 => CSA_sum_5_23_0, in2 => CSA_carry_5_22_0, c_in => CSA_carry_3_22_0, sum => CSA_sum_6_23_0, c_out => CSA_carry_6_23_0);
FA_lbl_6_24_0: FA port map(in1 => CSA_sum_5_24_0, in2 => CSA_carry_5_23_0, c_in => CSA_carry_2_23_0, sum => CSA_sum_6_24_0, c_out => CSA_carry_6_24_0);
FA_lbl_6_25_0: FA port map(in1 => CSA_sum_5_25_0, in2 => CSA_carry_5_24_0, c_in => CSA_carry_3_24_0, sum => CSA_sum_6_25_0, c_out => CSA_carry_6_25_0);
FA_lbl_6_26_0: FA port map(in1 => CSA_sum_5_26_0, in2 => CSA_carry_5_25_0, c_in => CSA_carry_0_25_0, sum => CSA_sum_6_26_0, c_out => CSA_carry_6_26_0);
FA_lbl_6_27_0: FA port map(in1 => CSA_sum_5_27_0, in2 => CSA_carry_5_26_0, c_in => CSA_carry_4_26_0, sum => CSA_sum_6_27_0, c_out => CSA_carry_6_27_0);
FA_lbl_6_28_0: FA port map(in1 => CSA_sum_5_28_0, in2 => CSA_carry_5_27_0, c_in => CSA_carry_4_27_0, sum => CSA_sum_6_28_0, c_out => CSA_carry_6_28_0);
FA_lbl_6_29_0: FA port map(in1 => CSA_sum_5_29_0, in2 => CSA_carry_5_28_0, c_in => CSA_carry_4_28_0, sum => CSA_sum_6_29_0, c_out => CSA_carry_6_29_0);
FA_lbl_6_30_0: FA port map(in1 => CSA_sum_5_30_0, in2 => CSA_carry_5_29_0, c_in => CSA_carry_4_29_0, sum => CSA_sum_6_30_0, c_out => CSA_carry_6_30_0);
FA_lbl_6_31_0: FA port map(in1 => CSA_sum_5_31_0, in2 => CSA_carry_5_30_0, c_in => CSA_carry_4_30_0, sum => CSA_sum_6_31_0, c_out => CSA_carry_6_31_0);
FA_lbl_6_32_0: FA port map(in1 => CSA_sum_5_32_1, in2 => CSA_sum_5_32_0, c_in => CSA_carry_5_31_0, sum => CSA_sum_6_32_0, c_out => CSA_carry_6_32_0);
FA_lbl_6_33_0: FA port map(in1 => CSA_sum_5_33_0, in2 => CSA_carry_5_32_1, c_in => CSA_carry_5_32_0, sum => CSA_sum_6_33_0, c_out => CSA_carry_6_33_0);
FA_lbl_6_34_0: FA port map(in1 => CSA_sum_5_34_0, in2 => CSA_carry_5_33_0, c_in => CSA_carry_4_33_0, sum => CSA_sum_6_34_0, c_out => CSA_carry_6_34_0);
FA_lbl_6_35_0: FA port map(in1 => CSA_sum_5_35_0, in2 => CSA_carry_5_34_0, c_in => CSA_carry_4_34_0, sum => CSA_sum_6_35_0, c_out => CSA_carry_6_35_0);
FA_lbl_6_36_0: FA port map(in1 => CSA_sum_5_36_0, in2 => CSA_carry_5_35_0, c_in => CSA_carry_4_35_0, sum => CSA_sum_6_36_0, c_out => CSA_carry_6_36_0);
FA_lbl_6_37_0: FA port map(in1 => CSA_sum_5_37_0, in2 => CSA_carry_5_36_0, c_in => CSA_carry_3_36_1, sum => CSA_sum_6_37_0, c_out => CSA_carry_6_37_0);
FA_lbl_6_39_0: FA port map(in1 => CSA_sum_5_39_0, in2 => CSA_carry_5_38_0, c_in => CSA_carry_4_38_0, sum => CSA_sum_6_39_0, c_out => CSA_carry_6_39_0);
FA_lbl_6_40_0: FA port map(in1 => CSA_sum_5_40_0, in2 => CSA_carry_5_39_0, c_in => CSA_carry_4_39_0, sum => CSA_sum_6_40_0, c_out => CSA_carry_6_40_0);
FA_lbl_6_41_0: FA port map(in1 => CSA_sum_5_41_0, in2 => CSA_carry_5_40_0, c_in => CSA_carry_4_40_0, sum => CSA_sum_6_41_0, c_out => CSA_carry_6_41_0);
FA_lbl_6_42_0: FA port map(in1 => CSA_sum_5_42_0, in2 => CSA_carry_5_41_0, c_in => CSA_carry_4_41_0, sum => CSA_sum_6_42_0, c_out => CSA_carry_6_42_0);
FA_lbl_6_43_0: FA port map(in1 => CSA_sum_5_43_0, in2 => CSA_carry_5_42_0, c_in => CSA_carry_3_42_0, sum => CSA_sum_6_43_0, c_out => CSA_carry_6_43_0);
FA_lbl_6_44_0: FA port map(in1 => CSA_sum_5_44_0, in2 => CSA_carry_5_43_0, c_in => CSA_carry_0_43_0, sum => CSA_sum_6_44_0, c_out => CSA_carry_6_44_0);
FA_lbl_6_45_0: FA port map(in1 => CSA_sum_5_45_0, in2 => CSA_carry_5_44_0, c_in => CSA_carry_1_44_0, sum => CSA_sum_6_45_0, c_out => CSA_carry_6_45_0);
FA_lbl_6_46_0: FA port map(in1 => CSA_sum_5_46_0, in2 => CSA_carry_5_45_0, c_in => CSA_carry_2_45_0, sum => CSA_sum_6_46_0, c_out => CSA_carry_6_46_0);
FA_lbl_6_47_0: FA port map(in1 => CSA_carry_5_46_0, in2 => CSA_sum_4_47_0, c_in => CSA_carry_4_46_0, sum => CSA_sum_6_47_0, c_out => CSA_carry_6_47_0);
FA_lbl_7_9_0: FA port map(in1 => CSA_carry_6_8_0, in2 => CSA_sum_3_9_0, c_in => CSA_carry_3_8_0, sum => CSA_sum_7_9_0, c_out => CSA_carry_7_9_0);
FA_lbl_7_33_0: FA port map(in1 => CSA_sum_6_33_0, in2 => CSA_carry_6_32_0, c_in => CSA_carry_4_32_0, sum => CSA_sum_7_33_0, c_out => CSA_carry_7_33_0);
FA_lbl_7_34_0: FA port map(in1 => CSA_sum_6_34_0, in2 => CSA_carry_6_33_0, c_in => CSA_carry_1_33_0, sum => CSA_sum_7_34_0, c_out => CSA_carry_7_34_0);
FA_lbl_7_35_0: FA port map(in1 => CSA_sum_6_35_0, in2 => CSA_carry_6_34_0, c_in => CSA_carry_0_34_0, sum => CSA_sum_7_35_0, c_out => CSA_carry_7_35_0);
FA_lbl_7_36_0: FA port map(in1 => CSA_sum_6_36_0, in2 => CSA_carry_6_35_0, c_in => CSA_carry_2_35_0, sum => CSA_sum_7_36_0, c_out => CSA_carry_7_36_0);
FA_lbl_7_37_0: FA port map(in1 => CSA_sum_6_37_0, in2 => CSA_carry_6_36_0, c_in => CSA_carry_3_36_0, sum => CSA_sum_7_37_0, c_out => CSA_carry_7_37_0);
FA_lbl_7_38_0: FA port map(in1 => CSA_carry_6_37_0, in2 => CSA_sum_5_38_0, c_in => CSA_carry_5_37_0, sum => CSA_sum_7_38_0, c_out => CSA_carry_7_38_0);
FA_lbl_8_10_0: FA port map(in1 => CSA_carry_7_9_0, in2 => CSA_sum_3_10_0, c_in => CSA_carry_3_9_0, sum => CSA_sum_8_10_0, c_out => CSA_carry_8_10_0);
FA_lbl_9_11_0: FA port map(in1 => CSA_carry_8_10_0, in2 => CSA_sum_4_11_0, c_in => CSA_carry_0_10_0, sum => CSA_sum_9_11_0, c_out => CSA_carry_9_11_0);
FA_lbl_10_12_0: FA port map(in1 => CSA_carry_9_11_0, in2 => CSA_sum_4_12_0, c_in => CSA_carry_4_11_0, sum => CSA_sum_10_12_0, c_out => CSA_carry_10_12_0);
FA_lbl_11_13_0: FA port map(in1 => CSA_carry_10_12_0, in2 => CSA_sum_4_13_0, c_in => CSA_carry_4_12_0, sum => CSA_sum_11_13_0, c_out => CSA_carry_11_13_0);
FA_lbl_12_14_0: FA port map(in1 => CSA_carry_11_13_0, in2 => CSA_sum_4_14_0, c_in => CSA_carry_4_13_0, sum => CSA_sum_12_14_0, c_out => CSA_carry_12_14_0);
FA_lbl_13_15_0: FA port map(in1 => CSA_carry_12_14_0, in2 => CSA_sum_4_15_0, c_in => CSA_carry_4_14_0, sum => CSA_sum_13_15_0, c_out => CSA_carry_13_15_0);
FA_lbl_14_16_0: FA port map(in1 => CSA_carry_13_15_0, in2 => CSA_sum_5_16_0, c_in => CSA_carry_1_15_0, sum => CSA_sum_14_16_0, c_out => CSA_carry_14_16_0);
FA_lbl_15_17_0: FA port map(in1 => CSA_carry_14_16_0, in2 => CSA_sum_5_17_0, c_in => CSA_carry_5_16_0, sum => CSA_sum_15_17_0, c_out => CSA_carry_15_17_0);
FA_lbl_16_18_0: FA port map(in1 => CSA_carry_15_17_0, in2 => CSA_sum_5_18_0, c_in => CSA_carry_5_17_0, sum => CSA_sum_16_18_0, c_out => CSA_carry_16_18_0);
FA_lbl_17_19_0: FA port map(in1 => CSA_carry_16_18_0, in2 => CSA_sum_5_19_0, c_in => CSA_carry_5_18_0, sum => CSA_sum_17_19_0, c_out => CSA_carry_17_19_0);
FA_lbl_18_20_0: FA port map(in1 => CSA_carry_17_19_0, in2 => CSA_sum_5_20_0, c_in => CSA_carry_5_19_0, sum => CSA_sum_18_20_0, c_out => CSA_carry_18_20_0);
FA_lbl_19_21_0: FA port map(in1 => CSA_carry_18_20_0, in2 => CSA_sum_5_21_0, c_in => CSA_carry_5_20_0, sum => CSA_sum_19_21_0, c_out => CSA_carry_19_21_0);
FA_lbl_20_22_0: FA port map(in1 => CSA_carry_19_21_0, in2 => CSA_sum_5_22_0, c_in => CSA_carry_5_21_0, sum => CSA_sum_20_22_0, c_out => CSA_carry_20_22_0);
FA_lbl_21_23_0: FA port map(in1 => CSA_carry_20_22_0, in2 => CSA_sum_6_23_0, c_in => CSA_carry_1_22_0, sum => CSA_sum_21_23_0, c_out => CSA_carry_21_23_0);
FA_lbl_22_24_0: FA port map(in1 => CSA_carry_21_23_0, in2 => CSA_sum_6_24_0, c_in => CSA_carry_6_23_0, sum => CSA_sum_22_24_0, c_out => CSA_carry_22_24_0);
FA_lbl_23_25_0: FA port map(in1 => CSA_carry_22_24_0, in2 => CSA_sum_6_25_0, c_in => CSA_carry_6_24_0, sum => CSA_sum_23_25_0, c_out => CSA_carry_23_25_0);
FA_lbl_24_26_0: FA port map(in1 => CSA_carry_23_25_0, in2 => CSA_sum_6_26_0, c_in => CSA_carry_6_25_0, sum => CSA_sum_24_26_0, c_out => CSA_carry_24_26_0);
FA_lbl_25_27_0: FA port map(in1 => CSA_carry_24_26_0, in2 => CSA_sum_6_27_0, c_in => CSA_carry_6_26_0, sum => CSA_sum_25_27_0, c_out => CSA_carry_25_27_0);
FA_lbl_26_28_0: FA port map(in1 => CSA_carry_25_27_0, in2 => CSA_sum_6_28_0, c_in => CSA_carry_6_27_0, sum => CSA_sum_26_28_0, c_out => CSA_carry_26_28_0);
FA_lbl_27_29_0: FA port map(in1 => CSA_carry_26_28_0, in2 => CSA_sum_6_29_0, c_in => CSA_carry_6_28_0, sum => CSA_sum_27_29_0, c_out => CSA_carry_27_29_0);
FA_lbl_28_30_0: FA port map(in1 => CSA_carry_27_29_0, in2 => CSA_sum_6_30_0, c_in => CSA_carry_6_29_0, sum => CSA_sum_28_30_0, c_out => CSA_carry_28_30_0);
FA_lbl_29_31_0: FA port map(in1 => CSA_carry_28_30_0, in2 => CSA_sum_6_31_0, c_in => CSA_carry_6_30_0, sum => CSA_sum_29_31_0, c_out => CSA_carry_29_31_0);
FA_lbl_30_32_0: FA port map(in1 => CSA_carry_29_31_0, in2 => CSA_sum_6_32_0, c_in => CSA_carry_6_31_0, sum => CSA_sum_30_32_0, c_out => CSA_carry_30_32_0);
out1(0) <= b_and_a(0);
out2(0) <= '0';
out1(1) <= b_and_a(1);
out2(1) <= b_and_a(32);
out1(2) <= CSA_sum_0_2_0;
out2(2) <= '0';
out1(3) <= CSA_sum_1_3_0;
out2(3) <= '0';
out1(4) <= CSA_sum_2_4_0;
out2(4) <= '0';
out1(5) <= CSA_sum_3_5_0;
out2(5) <= '0';
out1(6) <= CSA_sum_4_6_0;
out2(6) <= '0';
out1(7) <= CSA_sum_5_7_0;
out2(7) <= '0';
out1(8) <= CSA_sum_6_8_0;
out2(8) <= '0';
out1(9) <= CSA_sum_7_9_0;
out2(9) <= '0';
out1(10) <= CSA_sum_8_10_0;
out2(10) <= '0';
out1(11) <= CSA_sum_9_11_0;
out2(11) <= '0';
out1(12) <= CSA_sum_10_12_0;
out2(12) <= '0';
out1(13) <= CSA_sum_11_13_0;
out2(13) <= '0';
out1(14) <= CSA_sum_12_14_0;
out2(14) <= '0';
out1(15) <= CSA_sum_13_15_0;
out2(15) <= '0';
out1(16) <= CSA_sum_14_16_0;
out2(16) <= '0';
out1(17) <= CSA_sum_15_17_0;
out2(17) <= '0';
out1(18) <= CSA_sum_16_18_0;
out2(18) <= '0';
out1(19) <= CSA_sum_17_19_0;
out2(19) <= '0';
out1(20) <= CSA_sum_18_20_0;
out2(20) <= '0';
out1(21) <= CSA_sum_19_21_0;
out2(21) <= '0';
out1(22) <= CSA_sum_20_22_0;
out2(22) <= '0';
out1(23) <= CSA_sum_21_23_0;
out2(23) <= '0';
out1(24) <= CSA_sum_22_24_0;
out2(24) <= '0';
out1(25) <= CSA_sum_23_25_0;
out2(25) <= '0';
out1(26) <= CSA_sum_24_26_0;
out2(26) <= '0';
out1(27) <= CSA_sum_25_27_0;
out2(27) <= '0';
out1(28) <= CSA_sum_26_28_0;
out2(28) <= '0';
out1(29) <= CSA_sum_27_29_0;
out2(29) <= '0';
out1(30) <= CSA_sum_28_30_0;
out2(30) <= '0';
out1(31) <= CSA_sum_29_31_0;
out2(31) <= '0';
out1(32) <= CSA_sum_30_32_0;
out2(32) <= '0';
out1(33) <= CSA_carry_30_32_0;
out2(33) <= CSA_sum_7_33_0;
out1(34) <= CSA_sum_7_34_0;
out2(34) <= CSA_carry_7_33_0;
out1(35) <= CSA_sum_7_35_0;
out2(35) <= CSA_carry_7_34_0;
out1(36) <= CSA_sum_7_36_0;
out2(36) <= CSA_carry_7_35_0;
out1(37) <= CSA_sum_7_37_0;
out2(37) <= CSA_carry_7_36_0;
out1(38) <= CSA_sum_7_38_0;
out2(38) <= CSA_carry_7_37_0;
out1(39) <= CSA_carry_7_38_0;
out2(39) <= CSA_sum_6_39_0;
out1(40) <= CSA_sum_6_40_0;
out2(40) <= CSA_carry_6_39_0;
out1(41) <= CSA_sum_6_41_0;
out2(41) <= CSA_carry_6_40_0;
out1(42) <= CSA_sum_6_42_0;
out2(42) <= CSA_carry_6_41_0;
out1(43) <= CSA_sum_6_43_0;
out2(43) <= CSA_carry_6_42_0;
out1(44) <= CSA_sum_6_44_0;
out2(44) <= CSA_carry_6_43_0;
out1(45) <= CSA_sum_6_45_0;
out2(45) <= CSA_carry_6_44_0;
out1(46) <= CSA_sum_6_46_0;
out2(46) <= CSA_carry_6_45_0;
out1(47) <= CSA_sum_6_47_0;
out2(47) <= CSA_carry_6_46_0;
out1(48) <= CSA_carry_6_47_0;
out2(48) <= CSA_sum_5_48_0;
out1(49) <= CSA_sum_5_49_0;
out2(49) <= CSA_carry_5_48_0;
out1(50) <= CSA_sum_5_50_0;
out2(50) <= CSA_carry_5_49_0;
out1(51) <= CSA_sum_5_51_0;
out2(51) <= CSA_carry_5_50_0;
out1(52) <= CSA_sum_5_52_0;
out2(52) <= CSA_carry_5_51_0;
out1(53) <= CSA_sum_5_53_0;
out2(53) <= CSA_carry_5_52_0;
out1(54) <= CSA_carry_5_53_0;
out2(54) <= CSA_sum_4_54_0;
out1(55) <= CSA_sum_4_55_0;
out2(55) <= CSA_carry_4_54_0;
out1(56) <= CSA_sum_4_56_0;
out2(56) <= CSA_carry_4_55_0;
out1(57) <= CSA_sum_4_57_0;
out2(57) <= CSA_carry_4_56_0;
out1(58) <= CSA_carry_4_57_0;
out2(58) <= CSA_sum_3_58_0;
out1(59) <= CSA_sum_3_59_0;
out2(59) <= CSA_carry_3_58_0;
out1(60) <= CSA_carry_3_59_0;
out2(60) <= CSA_sum_2_60_0;
out1(61) <= CSA_carry_2_60_0;
out2(61) <= CSA_sum_1_61_0;
out1(62) <= CSA_carry_1_61_0;
out2(62) <= b_and_a(1023);
 end;